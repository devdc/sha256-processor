//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: Post-PnR Simulation Model file
//Tool Version: V1.9.9.03 (64-bit)
//Created Time: Tue Jun  3 12:23:31 2025

`timescale 100 ps/100 ps
module top_wrapper_tang9k(
	clk,
	rst,
	uart_rx,
	uart_tx,
	led0
);
input clk;
input rst;
input uart_rx;
output uart_tx;
output led0;
wire GND;
wire VCC;
wire clk;
wire led0;
wire rst;
wire uart_rx;
wire uart_tx;
wire \top/n568_23 ;
wire \top/tx_data_4_15 ;
wire \top/n636_5 ;
wire \top/data_in_7_6 ;
wire \top/send_index_6_7 ;
wire \top/n568_25 ;
wire \top/n585_15 ;
wire \top/n584_14 ;
wire \top/n582_14 ;
wire \top/n581_14 ;
wire \top/n580_14 ;
wire \top/n579_15 ;
wire \top/n567_20 ;
wire \top/n522_5 ;
wire \top/n523_5 ;
wire \top/n523_6 ;
wire \top/n525_4 ;
wire \top/n586_10 ;
wire \top/state_0_9 ;
wire \top/send_index_6_8 ;
wire \top/n568_26 ;
wire \top/n568_27 ;
wire \top/n568_28 ;
wire \top/n583_15 ;
wire \top/n580_15 ;
wire \top/n522_6 ;
wire \top/n522_7 ;
wire \top/n522_8 ;
wire \top/n522_9 ;
wire \top/n523_7 ;
wire \top/n523_8 ;
wire \top/n523_9 ;
wire \top/n523_10 ;
wire \top/n523_11 ;
wire \top/n523_12 ;
wire \top/n523_13 ;
wire \top/n523_14 ;
wire \top/n525_5 ;
wire \top/n525_6 ;
wire \top/n525_7 ;
wire \top/n525_8 ;
wire \top/n568_29 ;
wire \top/n568_30 ;
wire \top/n568_31 ;
wire \top/n568_32 ;
wire \top/n568_33 ;
wire \top/n522_10 ;
wire \top/n522_11 ;
wire \top/n522_12 ;
wire \top/n522_13 ;
wire \top/n522_14 ;
wire \top/n522_16 ;
wire \top/n522_17 ;
wire \top/n522_18 ;
wire \top/n522_19 ;
wire \top/n522_20 ;
wire \top/n522_21 ;
wire \top/n522_22 ;
wire \top/n522_23 ;
wire \top/n522_24 ;
wire \top/n522_25 ;
wire \top/n523_15 ;
wire \top/n523_16 ;
wire \top/n523_17 ;
wire \top/n523_18 ;
wire \top/n523_19 ;
wire \top/n523_20 ;
wire \top/n523_21 ;
wire \top/n523_22 ;
wire \top/n523_23 ;
wire \top/n523_24 ;
wire \top/n523_25 ;
wire \top/n523_26 ;
wire \top/n523_27 ;
wire \top/n523_28 ;
wire \top/n523_29 ;
wire \top/n523_30 ;
wire \top/n523_31 ;
wire \top/n523_32 ;
wire \top/n523_33 ;
wire \top/n523_34 ;
wire \top/n523_35 ;
wire \top/n523_36 ;
wire \top/n523_37 ;
wire \top/n523_38 ;
wire \top/n523_39 ;
wire \top/n523_40 ;
wire \top/n523_41 ;
wire \top/n523_42 ;
wire \top/n523_43 ;
wire \top/n523_44 ;
wire \top/n523_45 ;
wire \top/n523_46 ;
wire \top/n525_9 ;
wire \top/n525_10 ;
wire \top/n525_11 ;
wire \top/n525_12 ;
wire \top/n525_13 ;
wire \top/n525_14 ;
wire \top/n525_15 ;
wire \top/n525_16 ;
wire \top/n525_17 ;
wire \top/n525_18 ;
wire \top/n525_19 ;
wire \top/n525_20 ;
wire \top/n525_21 ;
wire \top/n525_22 ;
wire \top/n525_23 ;
wire \top/n525_24 ;
wire \top/n568_34 ;
wire \top/n522_26 ;
wire \top/n522_27 ;
wire \top/n522_28 ;
wire \top/n522_29 ;
wire \top/n522_30 ;
wire \top/n522_31 ;
wire \top/n522_32 ;
wire \top/n522_33 ;
wire \top/n522_34 ;
wire \top/n522_35 ;
wire \top/n522_36 ;
wire \top/n522_37 ;
wire \top/n522_38 ;
wire \top/n522_39 ;
wire \top/n522_40 ;
wire \top/n522_41 ;
wire \top/n522_42 ;
wire \top/n522_43 ;
wire \top/n522_44 ;
wire \top/n522_45 ;
wire \top/n522_46 ;
wire \top/n522_47 ;
wire \top/n522_48 ;
wire \top/n522_49 ;
wire \top/n522_50 ;
wire \top/n522_51 ;
wire \top/n522_52 ;
wire \top/n522_53 ;
wire \top/n522_54 ;
wire \top/n522_56 ;
wire \top/n522_57 ;
wire \top/n522_59 ;
wire \top/n522_60 ;
wire \top/n522_61 ;
wire \top/n522_62 ;
wire \top/n522_63 ;
wire \top/n522_64 ;
wire \top/n522_65 ;
wire \top/n522_66 ;
wire \top/n522_67 ;
wire \top/n522_68 ;
wire \top/n522_69 ;
wire \top/n522_70 ;
wire \top/n522_71 ;
wire \top/n522_72 ;
wire \top/n522_73 ;
wire \top/n523_47 ;
wire \top/n523_48 ;
wire \top/n523_49 ;
wire \top/n523_50 ;
wire \top/n523_52 ;
wire \top/n523_53 ;
wire \top/n523_54 ;
wire \top/n523_55 ;
wire \top/n523_56 ;
wire \top/n523_57 ;
wire \top/n523_59 ;
wire \top/n523_60 ;
wire \top/n523_61 ;
wire \top/n523_62 ;
wire \top/n523_63 ;
wire \top/n523_64 ;
wire \top/n523_65 ;
wire \top/n523_66 ;
wire \top/n523_67 ;
wire \top/n523_68 ;
wire \top/n523_69 ;
wire \top/n523_70 ;
wire \top/n523_71 ;
wire \top/n523_72 ;
wire \top/n523_73 ;
wire \top/n523_74 ;
wire \top/n523_75 ;
wire \top/n523_76 ;
wire \top/n523_77 ;
wire \top/n523_78 ;
wire \top/n523_79 ;
wire \top/n523_80 ;
wire \top/n523_81 ;
wire \top/n523_82 ;
wire \top/n523_83 ;
wire \top/n523_84 ;
wire \top/n523_85 ;
wire \top/n523_86 ;
wire \top/n523_87 ;
wire \top/n523_88 ;
wire \top/n523_89 ;
wire \top/n523_90 ;
wire \top/n523_91 ;
wire \top/n523_92 ;
wire \top/n523_93 ;
wire \top/n523_94 ;
wire \top/n523_95 ;
wire \top/n523_96 ;
wire \top/n523_97 ;
wire \top/n523_98 ;
wire \top/n523_99 ;
wire \top/n523_100 ;
wire \top/n523_102 ;
wire \top/n523_103 ;
wire \top/n523_104 ;
wire \top/n523_105 ;
wire \top/n523_106 ;
wire \top/n523_107 ;
wire \top/n523_108 ;
wire \top/n523_109 ;
wire \top/n523_110 ;
wire \top/n523_111 ;
wire \top/n523_112 ;
wire \top/n523_113 ;
wire \top/n523_114 ;
wire \top/n523_115 ;
wire \top/n523_116 ;
wire \top/n523_117 ;
wire \top/n523_118 ;
wire \top/n523_119 ;
wire \top/n525_25 ;
wire \top/n525_26 ;
wire \top/n525_27 ;
wire \top/n525_28 ;
wire \top/n525_29 ;
wire \top/n525_30 ;
wire \top/n525_31 ;
wire \top/n525_32 ;
wire \top/n525_33 ;
wire \top/n525_34 ;
wire \top/n525_35 ;
wire \top/n525_36 ;
wire \top/n525_37 ;
wire \top/n525_38 ;
wire \top/n525_39 ;
wire \top/n525_40 ;
wire \top/n525_41 ;
wire \top/n525_42 ;
wire \top/n525_43 ;
wire \top/n525_44 ;
wire \top/n525_45 ;
wire \top/n525_46 ;
wire \top/n525_47 ;
wire \top/n525_48 ;
wire \top/n525_49 ;
wire \top/n525_50 ;
wire \top/n525_51 ;
wire \top/n525_52 ;
wire \top/n525_53 ;
wire \top/n525_54 ;
wire \top/n525_55 ;
wire \top/n525_56 ;
wire \top/n525_57 ;
wire \top/n525_58 ;
wire \top/n525_59 ;
wire \top/n525_60 ;
wire \top/n525_61 ;
wire \top/n522_74 ;
wire \top/n522_75 ;
wire \top/n522_76 ;
wire \top/n522_77 ;
wire \top/n522_78 ;
wire \top/n522_79 ;
wire \top/n522_80 ;
wire \top/n522_81 ;
wire \top/n522_82 ;
wire \top/n522_83 ;
wire \top/n522_84 ;
wire \top/n522_85 ;
wire \top/n522_86 ;
wire \top/n523_120 ;
wire \top/n523_121 ;
wire \top/n523_122 ;
wire \top/n523_123 ;
wire \top/n523_124 ;
wire \top/n523_125 ;
wire \top/n523_126 ;
wire \top/n523_127 ;
wire \top/n523_128 ;
wire \top/n523_129 ;
wire \top/n523_130 ;
wire \top/n523_131 ;
wire \top/n523_132 ;
wire \top/n523_133 ;
wire \top/n523_134 ;
wire \top/n523_135 ;
wire \top/n523_136 ;
wire \top/n523_137 ;
wire \top/n523_138 ;
wire \top/n523_139 ;
wire \top/n523_140 ;
wire \top/n523_141 ;
wire \top/n523_142 ;
wire \top/n523_143 ;
wire \top/n523_144 ;
wire \top/n523_145 ;
wire \top/n525_62 ;
wire \top/n525_63 ;
wire \top/n525_64 ;
wire \top/n525_65 ;
wire \top/n525_66 ;
wire \top/n525_67 ;
wire \top/n525_68 ;
wire \top/n525_69 ;
wire \top/n525_70 ;
wire \top/n525_71 ;
wire \top/n525_72 ;
wire \top/n525_73 ;
wire \top/n525_74 ;
wire \top/n525_75 ;
wire \top/n524_5 ;
wire \top/n523_147 ;
wire \top/n570_11 ;
wire \top/tx_data_4_19 ;
wire \top/tx_data_5_19 ;
wire \top/n603_10 ;
wire \top/n586_12 ;
wire \top/n523_149 ;
wire \top/n525_77 ;
wire \top/n522_90 ;
wire \top/n523_151 ;
wire \top/n522_92 ;
wire \top/n522_94 ;
wire \top/n523_153 ;
wire \top/n582_17 ;
wire \top/n583_17 ;
wire \top/n569_27 ;
wire \top/state_0_13 ;
wire \top/n522_96 ;
wire \top/data_valid ;
wire \top/data_last ;
wire \top/tx_start ;
wire \top/rx_valid_Z ;
wire \top/tx_busy_Z ;
wire [6:0] \top/send_index ;
wire [6:0] \top/tx_data ;
wire [7:0] \top/data_in ;
wire [2:0] \top/state ;
wire [7:0] \top/rx_data_Z ;
wire [2:0] \top/state_0 ;
wire [255:0] \top/hash_out ;
wire \top/uart_rx_inst/n200_12 ;
wire \top/uart_rx_inst/n191_9 ;
wire \top/uart_rx_inst/bit_cnt_3_8 ;
wire \top/uart_rx_inst/n139_4 ;
wire \top/uart_rx_inst/n217_11 ;
wire \top/uart_rx_inst/n215_11 ;
wire \top/uart_rx_inst/n214_11 ;
wire \top/uart_rx_inst/n211_11 ;
wire \top/uart_rx_inst/n208_11 ;
wire \top/uart_rx_inst/n207_11 ;
wire \top/uart_rx_inst/n206_11 ;
wire \top/uart_rx_inst/n205_11 ;
wire \top/uart_rx_inst/n204_11 ;
wire \top/uart_rx_inst/n203_11 ;
wire \top/uart_rx_inst/n202_11 ;
wire \top/uart_rx_inst/n229_12 ;
wire \top/uart_rx_inst/n228_11 ;
wire \top/uart_rx_inst/n227_11 ;
wire \top/uart_rx_inst/n226_11 ;
wire \top/uart_rx_inst/n225_11 ;
wire \top/uart_rx_inst/n224_11 ;
wire \top/uart_rx_inst/n223_11 ;
wire \top/uart_rx_inst/n222_11 ;
wire \top/uart_rx_inst/n221_11 ;
wire \top/uart_rx_inst/n220_11 ;
wire \top/uart_rx_inst/n219_11 ;
wire \top/uart_rx_inst/n218_12 ;
wire \top/uart_rx_inst/n19_6 ;
wire \top/uart_rx_inst/n18_6 ;
wire \top/uart_rx_inst/n16_6 ;
wire \top/uart_rx_inst/n15_6 ;
wire \top/uart_rx_inst/n191_10 ;
wire \top/uart_rx_inst/baud_cnt_15_9 ;
wire \top/uart_rx_inst/state_0_10 ;
wire \top/uart_rx_inst/n214_12 ;
wire \top/uart_rx_inst/n211_12 ;
wire \top/uart_rx_inst/n208_12 ;
wire \top/uart_rx_inst/n206_12 ;
wire \top/uart_rx_inst/n204_12 ;
wire \top/uart_rx_inst/n203_12 ;
wire \top/uart_rx_inst/n226_12 ;
wire \top/uart_rx_inst/n18_7 ;
wire \top/uart_rx_inst/n15_7 ;
wire \top/uart_rx_inst/n191_11 ;
wire \top/uart_rx_inst/n191_12 ;
wire \top/uart_rx_inst/n191_13 ;
wire \top/uart_rx_inst/n191_14 ;
wire \top/uart_rx_inst/state_0_11 ;
wire \top/uart_rx_inst/rx_data_7_6 ;
wire \top/uart_rx_inst/shift_reg_7_10 ;
wire \top/uart_rx_inst/n217_14 ;
wire \top/uart_rx_inst/n22_8 ;
wire \top/uart_rx_inst/baud_cnt_8_9 ;
wire \top/uart_rx_inst/rx_d ;
wire \top/uart_rx_inst/rx_dd ;
wire \top/uart_rx_inst/rx_d_7 ;
wire \top/uart_rx_inst/n201_20 ;
wire [7:0] \top/uart_rx_inst/shift_reg ;
wire [3:0] \top/uart_rx_inst/bit_cnt ;
wire [15:0] \top/uart_rx_inst/baud_cnt ;
wire [1:0] \top/uart_rx_inst/state ;
wire \top/uart_tx_inst/tx_5 ;
wire \top/uart_tx_inst/n113_11 ;
wire \top/uart_tx_inst/n112_11 ;
wire \top/uart_tx_inst/n110_11 ;
wire \top/uart_tx_inst/n109_11 ;
wire \top/uart_tx_inst/n108_11 ;
wire \top/uart_tx_inst/n107_11 ;
wire \top/uart_tx_inst/n106_11 ;
wire \top/uart_tx_inst/n104_11 ;
wire \top/uart_tx_inst/n103_11 ;
wire \top/uart_tx_inst/n102_11 ;
wire \top/uart_tx_inst/n101_11 ;
wire \top/uart_tx_inst/n100_11 ;
wire \top/uart_tx_inst/n99_11 ;
wire \top/uart_tx_inst/n98_13 ;
wire \top/uart_tx_inst/n126_10 ;
wire \top/uart_tx_inst/tx_6 ;
wire \top/uart_tx_inst/tx_7 ;
wire \top/uart_tx_inst/n111_12 ;
wire \top/uart_tx_inst/n107_12 ;
wire \top/uart_tx_inst/n106_12 ;
wire \top/uart_tx_inst/n105_12 ;
wire \top/uart_tx_inst/n102_12 ;
wire \top/uart_tx_inst/n100_12 ;
wire \top/uart_tx_inst/n99_12 ;
wire \top/uart_tx_inst/n129_11 ;
wire \top/uart_tx_inst/n125_11 ;
wire \top/uart_tx_inst/tx_8 ;
wire \top/uart_tx_inst/tx_9 ;
wire \top/uart_tx_inst/n103_14 ;
wire \top/uart_tx_inst/n105_14 ;
wire \top/uart_tx_inst/n109_14 ;
wire \top/uart_tx_inst/n111_14 ;
wire \top/uart_tx_inst/n81_8 ;
wire \top/uart_tx_inst/n124_12 ;
wire \top/uart_tx_inst/n125_13 ;
wire \top/uart_tx_inst/n127_12 ;
wire \top/uart_tx_inst/n128_13 ;
wire \top/uart_tx_inst/n129_13 ;
wire \top/uart_tx_inst/baud_cnt_15_10 ;
wire \top/uart_tx_inst/n98_15 ;
wire \top/uart_tx_inst/n123_10 ;
wire \top/uart_tx_inst/n122_10 ;
wire \top/uart_tx_inst/n121_10 ;
wire \top/uart_tx_inst/n120_10 ;
wire \top/uart_tx_inst/n119_10 ;
wire \top/uart_tx_inst/n118_10 ;
wire \top/uart_tx_inst/n117_10 ;
wire \top/uart_tx_inst/tx_busy_7 ;
wire \top/uart_tx_inst/tx_busy_9 ;
wire \top/uart_tx_inst/n80_7 ;
wire [1:0] \top/uart_tx_inst/state ;
wire [15:0] \top/uart_tx_inst/baud_cnt ;
wire [3:0] \top/uart_tx_inst/bit_index ;
wire [8:0] \top/uart_tx_inst/shift_reg ;
wire \top/processor/n7631_3 ;
wire \top/processor/n10817_14 ;
wire \top/processor/n10825_14 ;
wire \top/processor/n11265_12 ;
wire \top/processor/n11266_12 ;
wire \top/processor/n11267_12 ;
wire \top/processor/n11268_12 ;
wire \top/processor/n11269_12 ;
wire \top/processor/n11270_12 ;
wire \top/processor/n11271_12 ;
wire \top/processor/n11272_12 ;
wire \top/processor/n11273_12 ;
wire \top/processor/n11274_12 ;
wire \top/processor/n11275_12 ;
wire \top/processor/n11276_12 ;
wire \top/processor/n11277_12 ;
wire \top/processor/n11278_12 ;
wire \top/processor/n11279_12 ;
wire \top/processor/n11280_12 ;
wire \top/processor/n11281_12 ;
wire \top/processor/n11282_12 ;
wire \top/processor/n11283_12 ;
wire \top/processor/n11284_12 ;
wire \top/processor/n11285_12 ;
wire \top/processor/n11286_12 ;
wire \top/processor/n11287_12 ;
wire \top/processor/n11288_12 ;
wire \top/processor/n11289_12 ;
wire \top/processor/n11290_12 ;
wire \top/processor/n11291_12 ;
wire \top/processor/n11292_12 ;
wire \top/processor/n11293_12 ;
wire \top/processor/n11294_12 ;
wire \top/processor/n11295_12 ;
wire \top/processor/n11296_12 ;
wire \top/processor/n11297_12 ;
wire \top/processor/n11298_12 ;
wire \top/processor/n11299_12 ;
wire \top/processor/n11300_12 ;
wire \top/processor/n11301_12 ;
wire \top/processor/n11302_12 ;
wire \top/processor/n11303_12 ;
wire \top/processor/n11304_12 ;
wire \top/processor/n11305_12 ;
wire \top/processor/n11306_12 ;
wire \top/processor/n11307_12 ;
wire \top/processor/n11308_12 ;
wire \top/processor/n11309_12 ;
wire \top/processor/n11310_12 ;
wire \top/processor/n11311_12 ;
wire \top/processor/n11312_12 ;
wire \top/processor/n11313_12 ;
wire \top/processor/n11314_12 ;
wire \top/processor/n11315_12 ;
wire \top/processor/n11316_12 ;
wire \top/processor/n11317_12 ;
wire \top/processor/n11318_12 ;
wire \top/processor/n11319_12 ;
wire \top/processor/n11320_12 ;
wire \top/processor/n11321_12 ;
wire \top/processor/n11322_12 ;
wire \top/processor/n11323_12 ;
wire \top/processor/n11324_12 ;
wire \top/processor/n11325_12 ;
wire \top/processor/n11361_16 ;
wire \top/processor/n11363_16 ;
wire \top/processor/n11364_27 ;
wire \top/processor/n11362_17 ;
wire \top/processor/state_0_10 ;
wire \top/processor/byte_index_5_8 ;
wire \top/processor/core_start_8 ;
wire \top/processor/hash_state_255_7 ;
wire \top/processor/total_bits_63_8 ;
wire \top/processor/seen_last_8 ;
wire \top/processor/need_length_block_8 ;
wire \top/processor/pad_index_5_8 ;
wire \top/processor/block_buffer_503_8 ;
wire \top/processor/block_buffer_495_8 ;
wire \top/processor/block_buffer_487_8 ;
wire \top/processor/block_buffer_479_8 ;
wire \top/processor/block_buffer_471_8 ;
wire \top/processor/block_buffer_463_8 ;
wire \top/processor/block_buffer_455_8 ;
wire \top/processor/block_buffer_439_8 ;
wire \top/processor/block_buffer_431_8 ;
wire \top/processor/block_buffer_423_8 ;
wire \top/processor/block_buffer_415_8 ;
wire \top/processor/block_buffer_407_8 ;
wire \top/processor/block_buffer_399_8 ;
wire \top/processor/block_buffer_391_8 ;
wire \top/processor/block_buffer_375_8 ;
wire \top/processor/block_buffer_367_8 ;
wire \top/processor/block_buffer_359_8 ;
wire \top/processor/block_buffer_351_8 ;
wire \top/processor/block_buffer_343_8 ;
wire \top/processor/block_buffer_335_8 ;
wire \top/processor/block_buffer_327_8 ;
wire \top/processor/block_buffer_319_8 ;
wire \top/processor/block_buffer_311_8 ;
wire \top/processor/block_buffer_303_8 ;
wire \top/processor/block_buffer_295_8 ;
wire \top/processor/block_buffer_287_8 ;
wire \top/processor/block_buffer_279_8 ;
wire \top/processor/block_buffer_271_8 ;
wire \top/processor/block_buffer_263_8 ;
wire \top/processor/block_buffer_247_8 ;
wire \top/processor/block_buffer_239_8 ;
wire \top/processor/block_buffer_231_8 ;
wire \top/processor/block_buffer_223_8 ;
wire \top/processor/block_buffer_215_8 ;
wire \top/processor/block_buffer_207_8 ;
wire \top/processor/block_buffer_199_8 ;
wire \top/processor/block_buffer_191_8 ;
wire \top/processor/block_buffer_183_8 ;
wire \top/processor/block_buffer_175_8 ;
wire \top/processor/block_buffer_167_8 ;
wire \top/processor/block_buffer_159_8 ;
wire \top/processor/block_buffer_151_8 ;
wire \top/processor/block_buffer_143_8 ;
wire \top/processor/block_buffer_135_8 ;
wire \top/processor/block_buffer_127_8 ;
wire \top/processor/block_buffer_119_8 ;
wire \top/processor/block_buffer_111_8 ;
wire \top/processor/block_buffer_103_8 ;
wire \top/processor/block_buffer_95_8 ;
wire \top/processor/block_buffer_87_8 ;
wire \top/processor/block_buffer_79_8 ;
wire \top/processor/block_buffer_71_8 ;
wire \top/processor/block_buffer_63_8 ;
wire \top/processor/block_buffer_55_8 ;
wire \top/processor/block_buffer_47_8 ;
wire \top/processor/block_buffer_39_8 ;
wire \top/processor/block_buffer_31_8 ;
wire \top/processor/block_buffer_23_8 ;
wire \top/processor/block_buffer_15_8 ;
wire \top/processor/block_ready_8 ;
wire \top/processor/n11438_14 ;
wire \top/processor/n11437_14 ;
wire \top/processor/n11436_14 ;
wire \top/processor/n11435_14 ;
wire \top/processor/n11434_14 ;
wire \top/processor/n11433_14 ;
wire \top/processor/n11432_14 ;
wire \top/processor/n11431_14 ;
wire \top/processor/n11429_14 ;
wire \top/processor/n11428_14 ;
wire \top/processor/n11427_14 ;
wire \top/processor/n11426_14 ;
wire \top/processor/n11425_14 ;
wire \top/processor/n11424_14 ;
wire \top/processor/n11422_14 ;
wire \top/processor/n11421_14 ;
wire \top/processor/n11420_14 ;
wire \top/processor/n11419_14 ;
wire \top/processor/n11418_14 ;
wire \top/processor/n11417_14 ;
wire \top/processor/n11416_14 ;
wire \top/processor/n11415_14 ;
wire \top/processor/n11413_14 ;
wire \top/processor/n11412_14 ;
wire \top/processor/n11411_14 ;
wire \top/processor/n11410_14 ;
wire \top/processor/n11408_14 ;
wire \top/processor/n11407_14 ;
wire \top/processor/n11406_14 ;
wire \top/processor/n11405_14 ;
wire \top/processor/n11404_14 ;
wire \top/processor/n11403_14 ;
wire \top/processor/n11402_14 ;
wire \top/processor/n11401_14 ;
wire \top/processor/n11400_14 ;
wire \top/processor/n11399_14 ;
wire \top/processor/n11398_14 ;
wire \top/processor/n11397_14 ;
wire \top/processor/n11396_14 ;
wire \top/processor/n11395_14 ;
wire \top/processor/n11394_14 ;
wire \top/processor/n11393_14 ;
wire \top/processor/n11392_14 ;
wire \top/processor/n11391_14 ;
wire \top/processor/n11389_14 ;
wire \top/processor/n11388_14 ;
wire \top/processor/n11387_14 ;
wire \top/processor/n11386_14 ;
wire \top/processor/n11385_14 ;
wire \top/processor/n11384_14 ;
wire \top/processor/n11383_14 ;
wire \top/processor/n11382_14 ;
wire \top/processor/n11381_14 ;
wire \top/processor/n11380_14 ;
wire \top/processor/n11379_14 ;
wire \top/processor/n11378_14 ;
wire \top/processor/n11377_14 ;
wire \top/processor/n11376_14 ;
wire \top/processor/n11375_14 ;
wire \top/processor/n11374_14 ;
wire \top/processor/n11373_14 ;
wire \top/processor/n11372_14 ;
wire \top/processor/n11368_17 ;
wire \top/processor/n11366_17 ;
wire \top/processor/n10824_15 ;
wire \top/processor/n10823_15 ;
wire \top/processor/n10822_15 ;
wire \top/processor/n10821_15 ;
wire \top/processor/n10820_15 ;
wire \top/processor/n10819_15 ;
wire \top/processor/n10818_15 ;
wire \top/processor/n10815_15 ;
wire \top/processor/n10814_15 ;
wire \top/processor/n10811_15 ;
wire \top/processor/n10810_15 ;
wire \top/processor/n10809_15 ;
wire \top/processor/n10807_15 ;
wire \top/processor/n10804_15 ;
wire \top/processor/n10803_15 ;
wire \top/processor/n10800_15 ;
wire \top/processor/n10799_15 ;
wire \top/processor/n10798_15 ;
wire \top/processor/n10797_15 ;
wire \top/processor/n10796_15 ;
wire \top/processor/n10790_15 ;
wire \top/processor/n10787_15 ;
wire \top/processor/n10785_15 ;
wire \top/processor/n10782_15 ;
wire \top/processor/n10780_15 ;
wire \top/processor/n10778_15 ;
wire \top/processor/n10775_15 ;
wire \top/processor/n10774_15 ;
wire \top/processor/n10771_15 ;
wire \top/processor/n10766_15 ;
wire \top/processor/n10765_15 ;
wire \top/processor/n10764_15 ;
wire \top/processor/n10763_15 ;
wire \top/processor/n10762_15 ;
wire \top/processor/n10755_15 ;
wire \top/processor/n10754_15 ;
wire \top/processor/n10753_15 ;
wire \top/processor/n10752_15 ;
wire \top/processor/n10751_15 ;
wire \top/processor/n10748_15 ;
wire \top/processor/n10747_15 ;
wire \top/processor/n10746_15 ;
wire \top/processor/n10744_15 ;
wire \top/processor/n10743_15 ;
wire \top/processor/n10742_15 ;
wire \top/processor/n10740_15 ;
wire \top/processor/n10737_15 ;
wire \top/processor/n10735_15 ;
wire \top/processor/n10733_15 ;
wire \top/processor/n10732_15 ;
wire \top/processor/n10731_15 ;
wire \top/processor/n10730_15 ;
wire \top/processor/n10729_15 ;
wire \top/processor/n10726_15 ;
wire \top/processor/n10723_15 ;
wire \top/processor/n10722_15 ;
wire \top/processor/n10713_15 ;
wire \top/processor/n10712_15 ;
wire \top/processor/n10710_15 ;
wire \top/processor/n10709_15 ;
wire \top/processor/n10707_15 ;
wire \top/processor/n10705_15 ;
wire \top/processor/n10704_15 ;
wire \top/processor/n10700_15 ;
wire \top/processor/n10699_15 ;
wire \top/processor/n10698_15 ;
wire \top/processor/n10697_15 ;
wire \top/processor/n10695_15 ;
wire \top/processor/n10694_15 ;
wire \top/processor/n10693_15 ;
wire \top/processor/n10691_15 ;
wire \top/processor/n10689_15 ;
wire \top/processor/n10688_15 ;
wire \top/processor/n10686_15 ;
wire \top/processor/n10682_15 ;
wire \top/processor/n10681_15 ;
wire \top/processor/n10679_15 ;
wire \top/processor/n10677_15 ;
wire \top/processor/n10668_15 ;
wire \top/processor/n10667_15 ;
wire \top/processor/n10665_15 ;
wire \top/processor/n10663_15 ;
wire \top/processor/n10661_15 ;
wire \top/processor/n10660_15 ;
wire \top/processor/n10658_15 ;
wire \top/processor/n10656_15 ;
wire \top/processor/n10654_15 ;
wire \top/processor/n10653_15 ;
wire \top/processor/n10649_15 ;
wire \top/processor/n10646_15 ;
wire \top/processor/n10645_15 ;
wire \top/processor/n10640_15 ;
wire \top/processor/n10636_15 ;
wire \top/processor/n10633_15 ;
wire \top/processor/n10632_15 ;
wire \top/processor/n10631_15 ;
wire \top/processor/n10626_15 ;
wire \top/processor/n10625_15 ;
wire \top/processor/n10623_15 ;
wire \top/processor/n10621_15 ;
wire \top/processor/n10620_15 ;
wire \top/processor/n10619_15 ;
wire \top/processor/n10618_15 ;
wire \top/processor/n10616_15 ;
wire \top/processor/n10612_15 ;
wire \top/processor/n10610_15 ;
wire \top/processor/n10605_15 ;
wire \top/processor/n10604_15 ;
wire \top/processor/n10601_15 ;
wire \top/processor/n10598_15 ;
wire \top/processor/n10594_15 ;
wire \top/processor/n10589_15 ;
wire \top/processor/n10588_15 ;
wire \top/processor/n10585_15 ;
wire \top/processor/n10584_15 ;
wire \top/processor/n10581_15 ;
wire \top/processor/n10580_15 ;
wire \top/processor/n10575_15 ;
wire \top/processor/n10574_15 ;
wire \top/processor/n10572_15 ;
wire \top/processor/n10571_15 ;
wire \top/processor/n10570_15 ;
wire \top/processor/n10569_15 ;
wire \top/processor/n10568_15 ;
wire \top/processor/n10566_15 ;
wire \top/processor/n10564_15 ;
wire \top/processor/n10561_16 ;
wire \top/processor/n9789_16 ;
wire \top/processor/n8408_6 ;
wire \top/processor/n10816_16 ;
wire \top/processor/n10813_16 ;
wire \top/processor/n10812_16 ;
wire \top/processor/n10808_16 ;
wire \top/processor/n10806_16 ;
wire \top/processor/n10805_16 ;
wire \top/processor/n10802_16 ;
wire \top/processor/n10801_16 ;
wire \top/processor/n10795_16 ;
wire \top/processor/n10794_16 ;
wire \top/processor/n10793_16 ;
wire \top/processor/n10792_16 ;
wire \top/processor/n10791_16 ;
wire \top/processor/n10789_16 ;
wire \top/processor/n10788_16 ;
wire \top/processor/n10786_16 ;
wire \top/processor/n10784_16 ;
wire \top/processor/n10783_16 ;
wire \top/processor/n10781_16 ;
wire \top/processor/n10779_16 ;
wire \top/processor/n10777_16 ;
wire \top/processor/n10776_16 ;
wire \top/processor/n10773_16 ;
wire \top/processor/n10772_16 ;
wire \top/processor/n10770_16 ;
wire \top/processor/n10769_16 ;
wire \top/processor/n10768_16 ;
wire \top/processor/n10767_16 ;
wire \top/processor/n10761_16 ;
wire \top/processor/n10760_16 ;
wire \top/processor/n10759_16 ;
wire \top/processor/n10758_16 ;
wire \top/processor/n10757_16 ;
wire \top/processor/n10756_16 ;
wire \top/processor/n10750_16 ;
wire \top/processor/n10749_16 ;
wire \top/processor/n10745_16 ;
wire \top/processor/n10741_16 ;
wire \top/processor/n10739_16 ;
wire \top/processor/n10738_16 ;
wire \top/processor/n10736_16 ;
wire \top/processor/n10734_16 ;
wire \top/processor/n10728_16 ;
wire \top/processor/n10727_16 ;
wire \top/processor/n10725_16 ;
wire \top/processor/n10724_16 ;
wire \top/processor/n10721_16 ;
wire \top/processor/n10720_16 ;
wire \top/processor/n10719_16 ;
wire \top/processor/n10718_16 ;
wire \top/processor/n10717_16 ;
wire \top/processor/n10716_16 ;
wire \top/processor/n10715_16 ;
wire \top/processor/n10714_16 ;
wire \top/processor/n10711_16 ;
wire \top/processor/n10708_16 ;
wire \top/processor/n10706_16 ;
wire \top/processor/n10703_16 ;
wire \top/processor/n10702_16 ;
wire \top/processor/n10701_16 ;
wire \top/processor/n10696_16 ;
wire \top/processor/n10692_16 ;
wire \top/processor/n10690_16 ;
wire \top/processor/n10687_16 ;
wire \top/processor/n10685_16 ;
wire \top/processor/n10684_16 ;
wire \top/processor/n10683_16 ;
wire \top/processor/n10680_16 ;
wire \top/processor/n10678_16 ;
wire \top/processor/n10676_16 ;
wire \top/processor/n10675_16 ;
wire \top/processor/n10674_16 ;
wire \top/processor/n10673_16 ;
wire \top/processor/n10672_16 ;
wire \top/processor/n10671_16 ;
wire \top/processor/n10670_16 ;
wire \top/processor/n10669_16 ;
wire \top/processor/n10666_16 ;
wire \top/processor/n10664_16 ;
wire \top/processor/n10662_16 ;
wire \top/processor/n10659_16 ;
wire \top/processor/n10657_16 ;
wire \top/processor/n10655_16 ;
wire \top/processor/n10652_16 ;
wire \top/processor/n10651_16 ;
wire \top/processor/n10650_16 ;
wire \top/processor/n10648_16 ;
wire \top/processor/n10647_16 ;
wire \top/processor/n10644_16 ;
wire \top/processor/n10643_16 ;
wire \top/processor/n10642_16 ;
wire \top/processor/n10641_16 ;
wire \top/processor/n10639_16 ;
wire \top/processor/n10638_16 ;
wire \top/processor/n10637_16 ;
wire \top/processor/n10635_16 ;
wire \top/processor/n10634_16 ;
wire \top/processor/n10630_16 ;
wire \top/processor/n10629_16 ;
wire \top/processor/n10628_16 ;
wire \top/processor/n10627_16 ;
wire \top/processor/n10624_16 ;
wire \top/processor/n10622_16 ;
wire \top/processor/n10617_16 ;
wire \top/processor/n10615_16 ;
wire \top/processor/n10614_16 ;
wire \top/processor/n10613_16 ;
wire \top/processor/n10611_16 ;
wire \top/processor/n10609_16 ;
wire \top/processor/n10608_16 ;
wire \top/processor/n10607_16 ;
wire \top/processor/n10606_16 ;
wire \top/processor/n10603_16 ;
wire \top/processor/n10602_16 ;
wire \top/processor/n10600_16 ;
wire \top/processor/n10599_16 ;
wire \top/processor/n10597_16 ;
wire \top/processor/n10596_16 ;
wire \top/processor/n10595_16 ;
wire \top/processor/n10593_16 ;
wire \top/processor/n10592_16 ;
wire \top/processor/n10591_16 ;
wire \top/processor/n10590_16 ;
wire \top/processor/n10587_16 ;
wire \top/processor/n10586_16 ;
wire \top/processor/n10583_16 ;
wire \top/processor/n10582_16 ;
wire \top/processor/n10579_16 ;
wire \top/processor/n10578_16 ;
wire \top/processor/n10577_16 ;
wire \top/processor/n10576_16 ;
wire \top/processor/n10573_16 ;
wire \top/processor/n10567_16 ;
wire \top/processor/n10565_16 ;
wire \top/processor/n10563_16 ;
wire \top/processor/n10562_16 ;
wire \top/processor/n9790_11 ;
wire \top/processor/n10817_15 ;
wire \top/processor/n11265_13 ;
wire \top/processor/n11361_17 ;
wire \top/processor/n11364_28 ;
wire \top/processor/n11362_18 ;
wire \top/processor/state_1_9 ;
wire \top/processor/hash_state_255_8 ;
wire \top/processor/seen_last_9 ;
wire \top/processor/need_length_block_9 ;
wire \top/processor/need_length_block_10 ;
wire \top/processor/block_buffer_511_9 ;
wire \top/processor/block_buffer_511_10 ;
wire \top/processor/block_buffer_511_11 ;
wire \top/processor/block_buffer_503_9 ;
wire \top/processor/block_buffer_503_10 ;
wire \top/processor/block_buffer_503_11 ;
wire \top/processor/block_buffer_495_9 ;
wire \top/processor/block_buffer_495_11 ;
wire \top/processor/block_buffer_487_9 ;
wire \top/processor/block_buffer_487_10 ;
wire \top/processor/block_buffer_479_9 ;
wire \top/processor/block_buffer_479_10 ;
wire \top/processor/block_buffer_471_9 ;
wire \top/processor/block_buffer_471_10 ;
wire \top/processor/block_buffer_463_9 ;
wire \top/processor/block_buffer_463_10 ;
wire \top/processor/block_buffer_455_9 ;
wire \top/processor/block_buffer_455_10 ;
wire \top/processor/block_buffer_447_9 ;
wire \top/processor/block_buffer_439_9 ;
wire \top/processor/block_buffer_439_10 ;
wire \top/processor/block_buffer_439_11 ;
wire \top/processor/block_buffer_431_9 ;
wire \top/processor/block_buffer_431_10 ;
wire \top/processor/block_buffer_423_9 ;
wire \top/processor/block_buffer_423_10 ;
wire \top/processor/block_buffer_415_9 ;
wire \top/processor/block_buffer_415_10 ;
wire \top/processor/block_buffer_407_9 ;
wire \top/processor/block_buffer_407_10 ;
wire \top/processor/block_buffer_399_9 ;
wire \top/processor/block_buffer_399_10 ;
wire \top/processor/block_buffer_391_9 ;
wire \top/processor/block_buffer_391_10 ;
wire \top/processor/block_buffer_383_9 ;
wire \top/processor/block_buffer_375_9 ;
wire \top/processor/block_buffer_375_10 ;
wire \top/processor/block_buffer_367_9 ;
wire \top/processor/block_buffer_359_9 ;
wire \top/processor/block_buffer_351_9 ;
wire \top/processor/block_buffer_343_9 ;
wire \top/processor/block_buffer_335_9 ;
wire \top/processor/block_buffer_327_9 ;
wire \top/processor/block_buffer_319_9 ;
wire \top/processor/block_buffer_319_10 ;
wire \top/processor/block_buffer_319_11 ;
wire \top/processor/block_buffer_311_9 ;
wire \top/processor/block_buffer_303_9 ;
wire \top/processor/block_buffer_295_9 ;
wire \top/processor/block_buffer_287_9 ;
wire \top/processor/block_buffer_279_9 ;
wire \top/processor/block_buffer_271_9 ;
wire \top/processor/block_buffer_263_9 ;
wire \top/processor/block_buffer_255_9 ;
wire \top/processor/block_buffer_247_9 ;
wire \top/processor/block_buffer_247_10 ;
wire \top/processor/block_buffer_239_9 ;
wire \top/processor/block_buffer_231_9 ;
wire \top/processor/block_buffer_223_9 ;
wire \top/processor/block_buffer_215_9 ;
wire \top/processor/block_buffer_207_9 ;
wire \top/processor/block_buffer_199_9 ;
wire \top/processor/block_buffer_191_9 ;
wire \top/processor/block_buffer_191_10 ;
wire \top/processor/block_buffer_183_9 ;
wire \top/processor/block_buffer_175_9 ;
wire \top/processor/block_buffer_167_9 ;
wire \top/processor/block_buffer_159_9 ;
wire \top/processor/block_buffer_151_9 ;
wire \top/processor/block_buffer_143_9 ;
wire \top/processor/block_buffer_135_9 ;
wire \top/processor/block_buffer_127_9 ;
wire \top/processor/block_buffer_127_10 ;
wire \top/processor/block_buffer_119_9 ;
wire \top/processor/block_buffer_111_9 ;
wire \top/processor/block_buffer_103_9 ;
wire \top/processor/block_buffer_95_9 ;
wire \top/processor/block_buffer_87_9 ;
wire \top/processor/block_buffer_79_9 ;
wire \top/processor/block_buffer_71_9 ;
wire \top/processor/block_buffer_63_9 ;
wire \top/processor/block_buffer_63_10 ;
wire \top/processor/block_buffer_63_11 ;
wire \top/processor/block_buffer_55_9 ;
wire \top/processor/block_buffer_55_10 ;
wire \top/processor/block_buffer_47_9 ;
wire \top/processor/block_buffer_39_9 ;
wire \top/processor/block_buffer_31_9 ;
wire \top/processor/block_buffer_31_10 ;
wire \top/processor/block_buffer_23_9 ;
wire \top/processor/block_buffer_15_9 ;
wire \top/processor/block_buffer_7_9 ;
wire \top/processor/n11435_15 ;
wire \top/processor/n11434_15 ;
wire \top/processor/n11432_15 ;
wire \top/processor/n11431_15 ;
wire \top/processor/n11430_15 ;
wire \top/processor/n11428_15 ;
wire \top/processor/n11425_15 ;
wire \top/processor/n11423_15 ;
wire \top/processor/n11420_15 ;
wire \top/processor/n11418_15 ;
wire \top/processor/n11417_15 ;
wire \top/processor/n11416_15 ;
wire \top/processor/n11415_15 ;
wire \top/processor/n11414_15 ;
wire \top/processor/n11412_15 ;
wire \top/processor/n11411_15 ;
wire \top/processor/n11410_15 ;
wire \top/processor/n11409_15 ;
wire \top/processor/n11407_15 ;
wire \top/processor/n11405_15 ;
wire \top/processor/n11403_15 ;
wire \top/processor/n11400_15 ;
wire \top/processor/n11399_15 ;
wire \top/processor/n11398_15 ;
wire \top/processor/n11396_15 ;
wire \top/processor/n11395_15 ;
wire \top/processor/n11394_15 ;
wire \top/processor/n11392_15 ;
wire \top/processor/n11390_15 ;
wire \top/processor/n11388_15 ;
wire \top/processor/n11387_15 ;
wire \top/processor/n11385_15 ;
wire \top/processor/n11383_15 ;
wire \top/processor/n11382_15 ;
wire \top/processor/n11380_15 ;
wire \top/processor/n11377_15 ;
wire \top/processor/n11376_15 ;
wire \top/processor/n11375_15 ;
wire \top/processor/n11375_16 ;
wire \top/processor/n11374_17 ;
wire \top/processor/n11373_15 ;
wire \top/processor/n11373_16 ;
wire \top/processor/n11372_15 ;
wire \top/processor/n11372_16 ;
wire \top/processor/n11370_19 ;
wire \top/processor/n11362_19 ;
wire \top/processor/state_1_10 ;
wire \top/processor/block_buffer_511_12 ;
wire \top/processor/block_buffer_511_13 ;
wire \top/processor/block_buffer_447_10 ;
wire \top/processor/block_buffer_447_11 ;
wire \top/processor/block_buffer_439_12 ;
wire \top/processor/block_buffer_423_11 ;
wire \top/processor/block_buffer_407_11 ;
wire \top/processor/block_buffer_383_10 ;
wire \top/processor/block_buffer_383_11 ;
wire \top/processor/block_buffer_375_11 ;
wire \top/processor/block_buffer_255_10 ;
wire \top/processor/block_buffer_255_11 ;
wire \top/processor/block_buffer_247_11 ;
wire \top/processor/block_buffer_191_11 ;
wire \top/processor/block_buffer_127_11 ;
wire \top/processor/n11420_16 ;
wire \top/processor/n11405_16 ;
wire \top/processor/n11396_16 ;
wire \top/processor/n11392_16 ;
wire \top/processor/n11390_16 ;
wire \top/processor/n11385_16 ;
wire \top/processor/n11376_16 ;
wire \top/processor/n11374_18 ;
wire \top/processor/block_buffer_447_12 ;
wire \top/processor/n11410_17 ;
wire \top/processor/n11405_17 ;
wire \top/processor/n11379_17 ;
wire \top/processor/n11382_18 ;
wire \top/processor/n11409_17 ;
wire \top/processor/n9790_13 ;
wire \top/processor/block_buffer_399_13 ;
wire \top/processor/block_buffer_431_13 ;
wire \top/processor/n11390_18 ;
wire \top/processor/n11402_17 ;
wire \top/processor/n11427_17 ;
wire \top/processor/block_buffer_319_15 ;
wire \top/processor/block_buffer_263_12 ;
wire \top/processor/block_buffer_319_17 ;
wire \top/processor/n11374_20 ;
wire \top/processor/n11414_17 ;
wire \top/processor/n11410_19 ;
wire \top/processor/core_busy_8 ;
wire \top/processor/n9790_15 ;
wire \top/processor/n11424_17 ;
wire \top/processor/n11430_17 ;
wire \top/processor/n7631_8 ;
wire \top/processor/n11365_19 ;
wire \top/processor/n11367_19 ;
wire \top/processor/n11369_19 ;
wire \top/processor/n11370_21 ;
wire \top/processor/n7631_10 ;
wire \top/processor/n7631_12 ;
wire \top/processor/n11374_22 ;
wire \top/processor/block_buffer_495_13 ;
wire \top/processor/block_buffer_7_11 ;
wire \top/processor/block_buffer_255_13 ;
wire \top/processor/block_buffer_383_13 ;
wire \top/processor/block_buffer_447_14 ;
wire \top/processor/block_buffer_511_15 ;
wire \top/processor/n11378_17 ;
wire \top/processor/n11421_17 ;
wire \top/processor/n11423_17 ;
wire \top/processor/block_ready ;
wire \top/processor/core_use_init ;
wire \top/processor/core_busy ;
wire \top/processor/core_ready_prev ;
wire \top/processor/seen_last ;
wire \top/processor/need_length_block ;
wire \top/processor/core_start ;
wire \top/processor/core_ready ;
wire [5:0] \top/processor/byte_index ;
wire [511:0] \top/processor/core_block ;
wire [255:0] \top/processor/core_hash_init ;
wire [63:3] \top/processor/total_bits ;
wire [5:0] \top/processor/pad_index ;
wire [511:0] \top/processor/block_buffer ;
wire [255:0] \top/processor/core_hash_out ;
wire \top/processor/sha_core/n3494_148 ;
wire \top/processor/sha_core/n3866_101 ;
wire \top/processor/sha_core/n3607_133 ;
wire \top/processor/sha_core/n3608_133 ;
wire \top/processor/sha_core/n3609_133 ;
wire \top/processor/sha_core/n3610_133 ;
wire \top/processor/sha_core/n3611_133 ;
wire \top/processor/sha_core/n3612_133 ;
wire \top/processor/sha_core/n3613_133 ;
wire \top/processor/sha_core/n3614_133 ;
wire \top/processor/sha_core/n3615_133 ;
wire \top/processor/sha_core/n3616_133 ;
wire \top/processor/sha_core/n3617_133 ;
wire \top/processor/sha_core/n3618_133 ;
wire \top/processor/sha_core/n3619_133 ;
wire \top/processor/sha_core/n3620_133 ;
wire \top/processor/sha_core/n3621_133 ;
wire \top/processor/sha_core/n3494_135 ;
wire \top/processor/sha_core/n3866_103 ;
wire \top/processor/sha_core/n3622_133 ;
wire \top/processor/sha_core/n3623_133 ;
wire \top/processor/sha_core/n3624_133 ;
wire \top/processor/sha_core/n3625_133 ;
wire \top/processor/sha_core/n3626_133 ;
wire \top/processor/sha_core/n3627_133 ;
wire \top/processor/sha_core/n3628_133 ;
wire \top/processor/sha_core/n3629_133 ;
wire \top/processor/sha_core/n3630_133 ;
wire \top/processor/sha_core/n3631_133 ;
wire \top/processor/sha_core/n3632_133 ;
wire \top/processor/sha_core/n3633_133 ;
wire \top/processor/sha_core/n3634_133 ;
wire \top/processor/sha_core/n3635_133 ;
wire \top/processor/sha_core/n3636_133 ;
wire \top/processor/sha_core/n3637_133 ;
wire \top/processor/sha_core/n3638_133 ;
wire \top/processor/sha_core/n3494_137 ;
wire \top/processor/sha_core/n3866_105 ;
wire \top/processor/sha_core/n3494_139 ;
wire \top/processor/sha_core/n3866_107 ;
wire \top/processor/sha_core/n3607_135 ;
wire \top/processor/sha_core/n3608_135 ;
wire \top/processor/sha_core/n3609_135 ;
wire \top/processor/sha_core/n3610_135 ;
wire \top/processor/sha_core/n3611_135 ;
wire \top/processor/sha_core/n3612_135 ;
wire \top/processor/sha_core/n3613_135 ;
wire \top/processor/sha_core/n3614_135 ;
wire \top/processor/sha_core/n3615_135 ;
wire \top/processor/sha_core/n3616_135 ;
wire \top/processor/sha_core/n3617_135 ;
wire \top/processor/sha_core/n3494_141 ;
wire \top/processor/sha_core/n3866_109 ;
wire \top/processor/sha_core/n3618_135 ;
wire \top/processor/sha_core/n3619_135 ;
wire \top/processor/sha_core/n3620_135 ;
wire \top/processor/sha_core/n3621_135 ;
wire \top/processor/sha_core/n3622_135 ;
wire \top/processor/sha_core/n3623_135 ;
wire \top/processor/sha_core/n3624_135 ;
wire \top/processor/sha_core/n3625_135 ;
wire \top/processor/sha_core/n3626_135 ;
wire \top/processor/sha_core/n3627_135 ;
wire \top/processor/sha_core/n3628_135 ;
wire \top/processor/sha_core/n3629_135 ;
wire \top/processor/sha_core/n3630_135 ;
wire \top/processor/sha_core/n3631_135 ;
wire \top/processor/sha_core/n3632_135 ;
wire \top/processor/sha_core/n3633_135 ;
wire \top/processor/sha_core/n3634_135 ;
wire \top/processor/sha_core/n3635_135 ;
wire \top/processor/sha_core/n3636_135 ;
wire \top/processor/sha_core/n3637_135 ;
wire \top/processor/sha_core/n3494_143 ;
wire \top/processor/sha_core/n3866_111 ;
wire \top/processor/sha_core/n3638_135 ;
wire \top/processor/sha_core/n3495_133 ;
wire \top/processor/sha_core/n3867_101 ;
wire \top/processor/sha_core/n3607_137 ;
wire \top/processor/sha_core/n3608_137 ;
wire \top/processor/sha_core/n3609_137 ;
wire \top/processor/sha_core/n3610_137 ;
wire \top/processor/sha_core/n3611_137 ;
wire \top/processor/sha_core/n3612_137 ;
wire \top/processor/sha_core/n3613_137 ;
wire \top/processor/sha_core/n3495_135 ;
wire \top/processor/sha_core/n3867_103 ;
wire \top/processor/sha_core/n3614_137 ;
wire \top/processor/sha_core/n3615_137 ;
wire \top/processor/sha_core/n3616_137 ;
wire \top/processor/sha_core/n3617_137 ;
wire \top/processor/sha_core/n3618_137 ;
wire \top/processor/sha_core/n3619_137 ;
wire \top/processor/sha_core/n3620_137 ;
wire \top/processor/sha_core/n3621_137 ;
wire \top/processor/sha_core/n3622_137 ;
wire \top/processor/sha_core/n3623_137 ;
wire \top/processor/sha_core/n3624_137 ;
wire \top/processor/sha_core/n3625_137 ;
wire \top/processor/sha_core/n3626_137 ;
wire \top/processor/sha_core/n3627_137 ;
wire \top/processor/sha_core/n3628_137 ;
wire \top/processor/sha_core/n3629_137 ;
wire \top/processor/sha_core/n3630_137 ;
wire \top/processor/sha_core/n3631_137 ;
wire \top/processor/sha_core/n3632_137 ;
wire \top/processor/sha_core/n3633_137 ;
wire \top/processor/sha_core/n3495_137 ;
wire \top/processor/sha_core/n3867_105 ;
wire \top/processor/sha_core/n3634_137 ;
wire \top/processor/sha_core/n3635_137 ;
wire \top/processor/sha_core/n3636_137 ;
wire \top/processor/sha_core/n3637_137 ;
wire \top/processor/sha_core/n3638_137 ;
wire \top/processor/sha_core/n3495_139 ;
wire \top/processor/sha_core/n3867_107 ;
wire \top/processor/sha_core/n3488_133 ;
wire \top/processor/sha_core/n3860_101 ;
wire \top/processor/sha_core/n3607_139 ;
wire \top/processor/sha_core/n3608_139 ;
wire \top/processor/sha_core/n3609_139 ;
wire \top/processor/sha_core/n3495_141 ;
wire \top/processor/sha_core/n3867_109 ;
wire \top/processor/sha_core/n3610_139 ;
wire \top/processor/sha_core/n3611_139 ;
wire \top/processor/sha_core/n3612_139 ;
wire \top/processor/sha_core/n3613_139 ;
wire \top/processor/sha_core/n3614_139 ;
wire \top/processor/sha_core/n3615_139 ;
wire \top/processor/sha_core/n3616_139 ;
wire \top/processor/sha_core/n3617_139 ;
wire \top/processor/sha_core/n3618_139 ;
wire \top/processor/sha_core/n3619_139 ;
wire \top/processor/sha_core/n3620_139 ;
wire \top/processor/sha_core/n3621_139 ;
wire \top/processor/sha_core/n3622_139 ;
wire \top/processor/sha_core/n3623_139 ;
wire \top/processor/sha_core/n3624_139 ;
wire \top/processor/sha_core/n3625_139 ;
wire \top/processor/sha_core/n3626_139 ;
wire \top/processor/sha_core/n3627_139 ;
wire \top/processor/sha_core/n3628_139 ;
wire \top/processor/sha_core/n3629_139 ;
wire \top/processor/sha_core/n3495_143 ;
wire \top/processor/sha_core/n3867_111 ;
wire \top/processor/sha_core/n3630_139 ;
wire \top/processor/sha_core/n3631_139 ;
wire \top/processor/sha_core/n3632_139 ;
wire \top/processor/sha_core/n3633_139 ;
wire \top/processor/sha_core/n3634_139 ;
wire \top/processor/sha_core/n3635_139 ;
wire \top/processor/sha_core/n3636_139 ;
wire \top/processor/sha_core/n3637_139 ;
wire \top/processor/sha_core/n3638_139 ;
wire \top/processor/sha_core/n3495_145 ;
wire \top/processor/sha_core/n3867_113 ;
wire \top/processor/sha_core/n3495_147 ;
wire \top/processor/sha_core/n3867_115 ;
wire \top/processor/sha_core/n3607_141 ;
wire \top/processor/sha_core/n3608_141 ;
wire \top/processor/sha_core/n3609_141 ;
wire \top/processor/sha_core/n3610_141 ;
wire \top/processor/sha_core/n3611_141 ;
wire \top/processor/sha_core/n3612_141 ;
wire \top/processor/sha_core/n3613_141 ;
wire \top/processor/sha_core/n3614_141 ;
wire \top/processor/sha_core/n3615_141 ;
wire \top/processor/sha_core/n3616_141 ;
wire \top/processor/sha_core/n3617_141 ;
wire \top/processor/sha_core/n3618_141 ;
wire \top/processor/sha_core/n3619_141 ;
wire \top/processor/sha_core/n3620_141 ;
wire \top/processor/sha_core/n3621_141 ;
wire \top/processor/sha_core/n3622_141 ;
wire \top/processor/sha_core/n3623_141 ;
wire \top/processor/sha_core/n3624_141 ;
wire \top/processor/sha_core/n3625_141 ;
wire \top/processor/sha_core/n3496_133 ;
wire \top/processor/sha_core/n3868_101 ;
wire \top/processor/sha_core/n3626_141 ;
wire \top/processor/sha_core/n3627_141 ;
wire \top/processor/sha_core/n3628_141 ;
wire \top/processor/sha_core/n3629_141 ;
wire \top/processor/sha_core/n3630_141 ;
wire \top/processor/sha_core/n3631_141 ;
wire \top/processor/sha_core/n3632_141 ;
wire \top/processor/sha_core/n3633_141 ;
wire \top/processor/sha_core/n3634_141 ;
wire \top/processor/sha_core/n3635_141 ;
wire \top/processor/sha_core/n3636_141 ;
wire \top/processor/sha_core/n3637_141 ;
wire \top/processor/sha_core/n3638_141 ;
wire \top/processor/sha_core/n3496_135 ;
wire \top/processor/sha_core/n3868_103 ;
wire \top/processor/sha_core/n3496_137 ;
wire \top/processor/sha_core/n3868_105 ;
wire \top/processor/sha_core/n3607_143 ;
wire \top/processor/sha_core/n3608_143 ;
wire \top/processor/sha_core/n3609_143 ;
wire \top/processor/sha_core/n3610_143 ;
wire \top/processor/sha_core/n3611_143 ;
wire \top/processor/sha_core/n3612_143 ;
wire \top/processor/sha_core/n3613_143 ;
wire \top/processor/sha_core/n3614_143 ;
wire \top/processor/sha_core/n3615_143 ;
wire \top/processor/sha_core/n3616_143 ;
wire \top/processor/sha_core/n3617_143 ;
wire \top/processor/sha_core/n3618_143 ;
wire \top/processor/sha_core/n3619_143 ;
wire \top/processor/sha_core/n3620_143 ;
wire \top/processor/sha_core/n3621_143 ;
wire \top/processor/sha_core/n3496_139 ;
wire \top/processor/sha_core/n3868_107 ;
wire \top/processor/sha_core/n3622_143 ;
wire \top/processor/sha_core/n3623_143 ;
wire \top/processor/sha_core/n3624_143 ;
wire \top/processor/sha_core/n3625_143 ;
wire \top/processor/sha_core/n3626_143 ;
wire \top/processor/sha_core/n3627_143 ;
wire \top/processor/sha_core/n3628_143 ;
wire \top/processor/sha_core/n3629_143 ;
wire \top/processor/sha_core/n3630_143 ;
wire \top/processor/sha_core/n3631_143 ;
wire \top/processor/sha_core/n3632_143 ;
wire \top/processor/sha_core/n3633_143 ;
wire \top/processor/sha_core/n3634_143 ;
wire \top/processor/sha_core/n3635_143 ;
wire \top/processor/sha_core/n3636_143 ;
wire \top/processor/sha_core/n3637_143 ;
wire \top/processor/sha_core/n3638_143 ;
wire \top/processor/sha_core/n3496_141 ;
wire \top/processor/sha_core/n3868_109 ;
wire \top/processor/sha_core/n3496_143 ;
wire \top/processor/sha_core/n3868_111 ;
wire \top/processor/sha_core/n3488_135 ;
wire \top/processor/sha_core/n3860_103 ;
wire \top/processor/sha_core/n3607_145 ;
wire \top/processor/sha_core/n3608_145 ;
wire \top/processor/sha_core/n3609_145 ;
wire \top/processor/sha_core/n3610_145 ;
wire \top/processor/sha_core/n3611_145 ;
wire \top/processor/sha_core/n3612_145 ;
wire \top/processor/sha_core/n3613_145 ;
wire \top/processor/sha_core/n3614_145 ;
wire \top/processor/sha_core/n3615_145 ;
wire \top/processor/sha_core/n3616_145 ;
wire \top/processor/sha_core/n3617_145 ;
wire \top/processor/sha_core/n3496_145 ;
wire \top/processor/sha_core/n3868_113 ;
wire \top/processor/sha_core/n3618_145 ;
wire \top/processor/sha_core/n3619_145 ;
wire \top/processor/sha_core/n3620_145 ;
wire \top/processor/sha_core/n3621_145 ;
wire \top/processor/sha_core/n3622_145 ;
wire \top/processor/sha_core/n3623_145 ;
wire \top/processor/sha_core/n3624_145 ;
wire \top/processor/sha_core/n3625_145 ;
wire \top/processor/sha_core/n3626_145 ;
wire \top/processor/sha_core/n3627_145 ;
wire \top/processor/sha_core/n3628_145 ;
wire \top/processor/sha_core/n3629_145 ;
wire \top/processor/sha_core/n3630_145 ;
wire \top/processor/sha_core/n3631_145 ;
wire \top/processor/sha_core/n3632_145 ;
wire \top/processor/sha_core/n3633_145 ;
wire \top/processor/sha_core/n3634_145 ;
wire \top/processor/sha_core/n3635_145 ;
wire \top/processor/sha_core/n3636_145 ;
wire \top/processor/sha_core/n3637_145 ;
wire \top/processor/sha_core/n3496_147 ;
wire \top/processor/sha_core/n3868_115 ;
wire \top/processor/sha_core/n3638_145 ;
wire \top/processor/sha_core/n3497_133 ;
wire \top/processor/sha_core/n3869_101 ;
wire \top/processor/sha_core/n3607_147 ;
wire \top/processor/sha_core/n3608_147 ;
wire \top/processor/sha_core/n3609_147 ;
wire \top/processor/sha_core/n3610_147 ;
wire \top/processor/sha_core/n3611_147 ;
wire \top/processor/sha_core/n3612_147 ;
wire \top/processor/sha_core/n3613_147 ;
wire \top/processor/sha_core/n3497_135 ;
wire \top/processor/sha_core/n3869_103 ;
wire \top/processor/sha_core/n3614_147 ;
wire \top/processor/sha_core/n3615_147 ;
wire \top/processor/sha_core/n3616_147 ;
wire \top/processor/sha_core/n3617_147 ;
wire \top/processor/sha_core/n3618_147 ;
wire \top/processor/sha_core/n3619_147 ;
wire \top/processor/sha_core/n3620_147 ;
wire \top/processor/sha_core/n3621_147 ;
wire \top/processor/sha_core/n3622_147 ;
wire \top/processor/sha_core/n3623_147 ;
wire \top/processor/sha_core/n3624_147 ;
wire \top/processor/sha_core/n3625_147 ;
wire \top/processor/sha_core/n3626_147 ;
wire \top/processor/sha_core/n3627_147 ;
wire \top/processor/sha_core/n3628_147 ;
wire \top/processor/sha_core/n3629_147 ;
wire \top/processor/sha_core/n3630_147 ;
wire \top/processor/sha_core/n3631_147 ;
wire \top/processor/sha_core/n3632_147 ;
wire \top/processor/sha_core/n3633_147 ;
wire \top/processor/sha_core/n3497_137 ;
wire \top/processor/sha_core/n3869_105 ;
wire \top/processor/sha_core/n3634_147 ;
wire \top/processor/sha_core/n3635_147 ;
wire \top/processor/sha_core/n3636_147 ;
wire \top/processor/sha_core/n3637_147 ;
wire \top/processor/sha_core/n3638_147 ;
wire \top/processor/sha_core/n3497_139 ;
wire \top/processor/sha_core/n3869_107 ;
wire \top/processor/sha_core/n3497_141 ;
wire \top/processor/sha_core/n3869_109 ;
wire \top/processor/sha_core/n3497_143 ;
wire \top/processor/sha_core/n3869_111 ;
wire \top/processor/sha_core/n3497_145 ;
wire \top/processor/sha_core/n3869_113 ;
wire \top/processor/sha_core/n3497_147 ;
wire \top/processor/sha_core/n3869_115 ;
wire \top/processor/sha_core/n3488_137 ;
wire \top/processor/sha_core/n3860_105 ;
wire \top/processor/sha_core/n3498_133 ;
wire \top/processor/sha_core/n3870_101 ;
wire \top/processor/sha_core/n3498_135 ;
wire \top/processor/sha_core/n3870_103 ;
wire \top/processor/sha_core/n3498_137 ;
wire \top/processor/sha_core/n3870_105 ;
wire \top/processor/sha_core/n3498_139 ;
wire \top/processor/sha_core/n3870_107 ;
wire \top/processor/sha_core/n3498_141 ;
wire \top/processor/sha_core/n3870_109 ;
wire \top/processor/sha_core/n3498_143 ;
wire \top/processor/sha_core/n3870_111 ;
wire \top/processor/sha_core/n3498_145 ;
wire \top/processor/sha_core/n3870_113 ;
wire \top/processor/sha_core/n3498_147 ;
wire \top/processor/sha_core/n3870_115 ;
wire \top/processor/sha_core/n3499_133 ;
wire \top/processor/sha_core/n3871_101 ;
wire \top/processor/sha_core/n3499_135 ;
wire \top/processor/sha_core/n3871_103 ;
wire \top/processor/sha_core/n3489_133 ;
wire \top/processor/sha_core/n3861_101 ;
wire \top/processor/sha_core/n3499_137 ;
wire \top/processor/sha_core/n3871_105 ;
wire \top/processor/sha_core/n3499_139 ;
wire \top/processor/sha_core/n3871_107 ;
wire \top/processor/sha_core/n3499_141 ;
wire \top/processor/sha_core/n3871_109 ;
wire \top/processor/sha_core/n3499_143 ;
wire \top/processor/sha_core/n3871_111 ;
wire \top/processor/sha_core/n3499_145 ;
wire \top/processor/sha_core/n3871_113 ;
wire \top/processor/sha_core/n3499_147 ;
wire \top/processor/sha_core/n3871_115 ;
wire \top/processor/sha_core/n3500_133 ;
wire \top/processor/sha_core/n3872_101 ;
wire \top/processor/sha_core/n3500_135 ;
wire \top/processor/sha_core/n3872_103 ;
wire \top/processor/sha_core/n3500_137 ;
wire \top/processor/sha_core/n3872_105 ;
wire \top/processor/sha_core/n3500_139 ;
wire \top/processor/sha_core/n3872_107 ;
wire \top/processor/sha_core/n3489_135 ;
wire \top/processor/sha_core/n3861_103 ;
wire \top/processor/sha_core/n3488_139 ;
wire \top/processor/sha_core/n3860_107 ;
wire \top/processor/sha_core/n3500_141 ;
wire \top/processor/sha_core/n3872_109 ;
wire \top/processor/sha_core/n3500_143 ;
wire \top/processor/sha_core/n3872_111 ;
wire \top/processor/sha_core/n3500_145 ;
wire \top/processor/sha_core/n3872_113 ;
wire \top/processor/sha_core/n3500_147 ;
wire \top/processor/sha_core/n3872_115 ;
wire \top/processor/sha_core/n3501_133 ;
wire \top/processor/sha_core/n3873_101 ;
wire \top/processor/sha_core/n3501_135 ;
wire \top/processor/sha_core/n3873_103 ;
wire \top/processor/sha_core/n3501_137 ;
wire \top/processor/sha_core/n3873_105 ;
wire \top/processor/sha_core/n3501_139 ;
wire \top/processor/sha_core/n3873_107 ;
wire \top/processor/sha_core/n3501_141 ;
wire \top/processor/sha_core/n3873_109 ;
wire \top/processor/sha_core/n3501_143 ;
wire \top/processor/sha_core/n3873_111 ;
wire \top/processor/sha_core/n3489_137 ;
wire \top/processor/sha_core/n3861_105 ;
wire \top/processor/sha_core/n3501_145 ;
wire \top/processor/sha_core/n3873_113 ;
wire \top/processor/sha_core/n3501_147 ;
wire \top/processor/sha_core/n3873_115 ;
wire \top/processor/sha_core/n3502_133 ;
wire \top/processor/sha_core/n3874_101 ;
wire \top/processor/sha_core/n3502_135 ;
wire \top/processor/sha_core/n3874_103 ;
wire \top/processor/sha_core/n3502_137 ;
wire \top/processor/sha_core/n3874_105 ;
wire \top/processor/sha_core/n3502_139 ;
wire \top/processor/sha_core/n3874_107 ;
wire \top/processor/sha_core/n3502_141 ;
wire \top/processor/sha_core/n3874_109 ;
wire \top/processor/sha_core/n3502_143 ;
wire \top/processor/sha_core/n3874_111 ;
wire \top/processor/sha_core/n3502_145 ;
wire \top/processor/sha_core/n3874_113 ;
wire \top/processor/sha_core/n3502_147 ;
wire \top/processor/sha_core/n3874_115 ;
wire \top/processor/sha_core/n3489_139 ;
wire \top/processor/sha_core/n3861_107 ;
wire \top/processor/sha_core/n3503_133 ;
wire \top/processor/sha_core/n3875_101 ;
wire \top/processor/sha_core/n3503_135 ;
wire \top/processor/sha_core/n3875_103 ;
wire \top/processor/sha_core/n3503_137 ;
wire \top/processor/sha_core/n3875_105 ;
wire \top/processor/sha_core/n3503_139 ;
wire \top/processor/sha_core/n3875_107 ;
wire \top/processor/sha_core/n3503_141 ;
wire \top/processor/sha_core/n3875_109 ;
wire \top/processor/sha_core/n3503_143 ;
wire \top/processor/sha_core/n3875_111 ;
wire \top/processor/sha_core/n3503_145 ;
wire \top/processor/sha_core/n3875_113 ;
wire \top/processor/sha_core/n3503_147 ;
wire \top/processor/sha_core/n3875_115 ;
wire \top/processor/sha_core/n3504_133 ;
wire \top/processor/sha_core/n3876_101 ;
wire \top/processor/sha_core/n3504_135 ;
wire \top/processor/sha_core/n3876_103 ;
wire \top/processor/sha_core/n3489_141 ;
wire \top/processor/sha_core/n3861_109 ;
wire \top/processor/sha_core/n3504_137 ;
wire \top/processor/sha_core/n3876_105 ;
wire \top/processor/sha_core/n3504_139 ;
wire \top/processor/sha_core/n3876_107 ;
wire \top/processor/sha_core/n3504_141 ;
wire \top/processor/sha_core/n3876_109 ;
wire \top/processor/sha_core/n3504_143 ;
wire \top/processor/sha_core/n3876_111 ;
wire \top/processor/sha_core/n3504_145 ;
wire \top/processor/sha_core/n3876_113 ;
wire \top/processor/sha_core/n3504_147 ;
wire \top/processor/sha_core/n3876_115 ;
wire \top/processor/sha_core/n3505_133 ;
wire \top/processor/sha_core/n3877_101 ;
wire \top/processor/sha_core/n3505_135 ;
wire \top/processor/sha_core/n3877_103 ;
wire \top/processor/sha_core/n3505_137 ;
wire \top/processor/sha_core/n3877_105 ;
wire \top/processor/sha_core/n3505_139 ;
wire \top/processor/sha_core/n3877_107 ;
wire \top/processor/sha_core/n3489_143 ;
wire \top/processor/sha_core/n3861_111 ;
wire \top/processor/sha_core/n3505_141 ;
wire \top/processor/sha_core/n3877_109 ;
wire \top/processor/sha_core/n3505_143 ;
wire \top/processor/sha_core/n3877_111 ;
wire \top/processor/sha_core/n3505_145 ;
wire \top/processor/sha_core/n3877_113 ;
wire \top/processor/sha_core/n3505_147 ;
wire \top/processor/sha_core/n3877_115 ;
wire \top/processor/sha_core/n3506_133 ;
wire \top/processor/sha_core/n3878_101 ;
wire \top/processor/sha_core/n3506_135 ;
wire \top/processor/sha_core/n3878_103 ;
wire \top/processor/sha_core/n3506_137 ;
wire \top/processor/sha_core/n3878_105 ;
wire \top/processor/sha_core/n3506_139 ;
wire \top/processor/sha_core/n3878_107 ;
wire \top/processor/sha_core/n3506_141 ;
wire \top/processor/sha_core/n3878_109 ;
wire \top/processor/sha_core/n3506_143 ;
wire \top/processor/sha_core/n3878_111 ;
wire \top/processor/sha_core/n3489_145 ;
wire \top/processor/sha_core/n3861_113 ;
wire \top/processor/sha_core/n3506_145 ;
wire \top/processor/sha_core/n3878_113 ;
wire \top/processor/sha_core/n3506_147 ;
wire \top/processor/sha_core/n3878_115 ;
wire \top/processor/sha_core/n3507_133 ;
wire \top/processor/sha_core/n3879_101 ;
wire \top/processor/sha_core/n3507_135 ;
wire \top/processor/sha_core/n3879_103 ;
wire \top/processor/sha_core/n3507_137 ;
wire \top/processor/sha_core/n3879_105 ;
wire \top/processor/sha_core/n3507_139 ;
wire \top/processor/sha_core/n3879_107 ;
wire \top/processor/sha_core/n3507_141 ;
wire \top/processor/sha_core/n3879_109 ;
wire \top/processor/sha_core/n3507_143 ;
wire \top/processor/sha_core/n3879_111 ;
wire \top/processor/sha_core/n3507_145 ;
wire \top/processor/sha_core/n3879_113 ;
wire \top/processor/sha_core/n3507_147 ;
wire \top/processor/sha_core/n3879_115 ;
wire \top/processor/sha_core/n3489_147 ;
wire \top/processor/sha_core/n3861_115 ;
wire \top/processor/sha_core/n3508_133 ;
wire \top/processor/sha_core/n3880_101 ;
wire \top/processor/sha_core/n3508_135 ;
wire \top/processor/sha_core/n3880_103 ;
wire \top/processor/sha_core/n3508_137 ;
wire \top/processor/sha_core/n3880_105 ;
wire \top/processor/sha_core/n3508_139 ;
wire \top/processor/sha_core/n3880_107 ;
wire \top/processor/sha_core/n3508_141 ;
wire \top/processor/sha_core/n3880_109 ;
wire \top/processor/sha_core/n3508_143 ;
wire \top/processor/sha_core/n3880_111 ;
wire \top/processor/sha_core/n3508_145 ;
wire \top/processor/sha_core/n3880_113 ;
wire \top/processor/sha_core/n3508_147 ;
wire \top/processor/sha_core/n3880_115 ;
wire \top/processor/sha_core/n3509_133 ;
wire \top/processor/sha_core/n3881_101 ;
wire \top/processor/sha_core/n3509_135 ;
wire \top/processor/sha_core/n3881_103 ;
wire \top/processor/sha_core/n3490_133 ;
wire \top/processor/sha_core/n3862_101 ;
wire \top/processor/sha_core/n3509_137 ;
wire \top/processor/sha_core/n3881_105 ;
wire \top/processor/sha_core/n3509_139 ;
wire \top/processor/sha_core/n3881_107 ;
wire \top/processor/sha_core/n3509_141 ;
wire \top/processor/sha_core/n3881_109 ;
wire \top/processor/sha_core/n3509_143 ;
wire \top/processor/sha_core/n3881_111 ;
wire \top/processor/sha_core/n3509_145 ;
wire \top/processor/sha_core/n3881_113 ;
wire \top/processor/sha_core/n3509_147 ;
wire \top/processor/sha_core/n3881_115 ;
wire \top/processor/sha_core/n3510_133 ;
wire \top/processor/sha_core/n3882_101 ;
wire \top/processor/sha_core/n3510_135 ;
wire \top/processor/sha_core/n3882_103 ;
wire \top/processor/sha_core/n3510_137 ;
wire \top/processor/sha_core/n3882_105 ;
wire \top/processor/sha_core/n3510_139 ;
wire \top/processor/sha_core/n3882_107 ;
wire \top/processor/sha_core/n3490_135 ;
wire \top/processor/sha_core/n3862_103 ;
wire \top/processor/sha_core/n3510_141 ;
wire \top/processor/sha_core/n3882_109 ;
wire \top/processor/sha_core/n3510_143 ;
wire \top/processor/sha_core/n3882_111 ;
wire \top/processor/sha_core/n3510_145 ;
wire \top/processor/sha_core/n3882_113 ;
wire \top/processor/sha_core/n3510_147 ;
wire \top/processor/sha_core/n3882_115 ;
wire \top/processor/sha_core/n3511_133 ;
wire \top/processor/sha_core/n3883_101 ;
wire \top/processor/sha_core/n3511_135 ;
wire \top/processor/sha_core/n3883_103 ;
wire \top/processor/sha_core/n3511_137 ;
wire \top/processor/sha_core/n3883_105 ;
wire \top/processor/sha_core/n3511_139 ;
wire \top/processor/sha_core/n3883_107 ;
wire \top/processor/sha_core/n3511_141 ;
wire \top/processor/sha_core/n3883_109 ;
wire \top/processor/sha_core/n3511_143 ;
wire \top/processor/sha_core/n3883_111 ;
wire \top/processor/sha_core/n3490_137 ;
wire \top/processor/sha_core/n3862_105 ;
wire \top/processor/sha_core/n3511_145 ;
wire \top/processor/sha_core/n3883_113 ;
wire \top/processor/sha_core/n3511_147 ;
wire \top/processor/sha_core/n3883_115 ;
wire \top/processor/sha_core/n3512_133 ;
wire \top/processor/sha_core/n3884_101 ;
wire \top/processor/sha_core/n3512_135 ;
wire \top/processor/sha_core/n3884_103 ;
wire \top/processor/sha_core/n3512_137 ;
wire \top/processor/sha_core/n3884_105 ;
wire \top/processor/sha_core/n3512_139 ;
wire \top/processor/sha_core/n3884_107 ;
wire \top/processor/sha_core/n3512_141 ;
wire \top/processor/sha_core/n3884_109 ;
wire \top/processor/sha_core/n3512_143 ;
wire \top/processor/sha_core/n3884_111 ;
wire \top/processor/sha_core/n3512_145 ;
wire \top/processor/sha_core/n3884_113 ;
wire \top/processor/sha_core/n3512_147 ;
wire \top/processor/sha_core/n3884_115 ;
wire \top/processor/sha_core/n3490_139 ;
wire \top/processor/sha_core/n3862_107 ;
wire \top/processor/sha_core/n3488_141 ;
wire \top/processor/sha_core/n3860_109 ;
wire \top/processor/sha_core/n3513_133 ;
wire \top/processor/sha_core/n3885_101 ;
wire \top/processor/sha_core/n3513_135 ;
wire \top/processor/sha_core/n3885_103 ;
wire \top/processor/sha_core/n3513_137 ;
wire \top/processor/sha_core/n3885_105 ;
wire \top/processor/sha_core/n3513_139 ;
wire \top/processor/sha_core/n3885_107 ;
wire \top/processor/sha_core/n3513_141 ;
wire \top/processor/sha_core/n3885_109 ;
wire \top/processor/sha_core/n3513_143 ;
wire \top/processor/sha_core/n3885_111 ;
wire \top/processor/sha_core/n3513_145 ;
wire \top/processor/sha_core/n3885_113 ;
wire \top/processor/sha_core/n3513_147 ;
wire \top/processor/sha_core/n3885_115 ;
wire \top/processor/sha_core/n3514_133 ;
wire \top/processor/sha_core/n3886_101 ;
wire \top/processor/sha_core/n3514_135 ;
wire \top/processor/sha_core/n3886_103 ;
wire \top/processor/sha_core/n3490_141 ;
wire \top/processor/sha_core/n3862_109 ;
wire \top/processor/sha_core/n3514_137 ;
wire \top/processor/sha_core/n3886_105 ;
wire \top/processor/sha_core/n3514_139 ;
wire \top/processor/sha_core/n3886_107 ;
wire \top/processor/sha_core/n3514_141 ;
wire \top/processor/sha_core/n3886_109 ;
wire \top/processor/sha_core/n3514_143 ;
wire \top/processor/sha_core/n3886_111 ;
wire \top/processor/sha_core/n3514_145 ;
wire \top/processor/sha_core/n3886_113 ;
wire \top/processor/sha_core/n3514_147 ;
wire \top/processor/sha_core/n3886_115 ;
wire \top/processor/sha_core/n3515_133 ;
wire \top/processor/sha_core/n3887_101 ;
wire \top/processor/sha_core/n3515_135 ;
wire \top/processor/sha_core/n3887_103 ;
wire \top/processor/sha_core/n3515_137 ;
wire \top/processor/sha_core/n3887_105 ;
wire \top/processor/sha_core/n3515_139 ;
wire \top/processor/sha_core/n3887_107 ;
wire \top/processor/sha_core/n3490_143 ;
wire \top/processor/sha_core/n3862_111 ;
wire \top/processor/sha_core/n3515_141 ;
wire \top/processor/sha_core/n3887_109 ;
wire \top/processor/sha_core/n3515_143 ;
wire \top/processor/sha_core/n3887_111 ;
wire \top/processor/sha_core/n3515_145 ;
wire \top/processor/sha_core/n3887_113 ;
wire \top/processor/sha_core/n3515_147 ;
wire \top/processor/sha_core/n3887_115 ;
wire \top/processor/sha_core/n3516_133 ;
wire \top/processor/sha_core/n3888_101 ;
wire \top/processor/sha_core/n3516_135 ;
wire \top/processor/sha_core/n3888_103 ;
wire \top/processor/sha_core/n3516_137 ;
wire \top/processor/sha_core/n3888_105 ;
wire \top/processor/sha_core/n3516_139 ;
wire \top/processor/sha_core/n3888_107 ;
wire \top/processor/sha_core/n3516_141 ;
wire \top/processor/sha_core/n3888_109 ;
wire \top/processor/sha_core/n3516_143 ;
wire \top/processor/sha_core/n3888_111 ;
wire \top/processor/sha_core/n3490_145 ;
wire \top/processor/sha_core/n3862_113 ;
wire \top/processor/sha_core/n3516_145 ;
wire \top/processor/sha_core/n3888_113 ;
wire \top/processor/sha_core/n3516_147 ;
wire \top/processor/sha_core/n3888_115 ;
wire \top/processor/sha_core/n3517_133 ;
wire \top/processor/sha_core/n3889_101 ;
wire \top/processor/sha_core/n3517_135 ;
wire \top/processor/sha_core/n3889_103 ;
wire \top/processor/sha_core/n3517_137 ;
wire \top/processor/sha_core/n3889_105 ;
wire \top/processor/sha_core/n3517_139 ;
wire \top/processor/sha_core/n3889_107 ;
wire \top/processor/sha_core/n3517_141 ;
wire \top/processor/sha_core/n3889_109 ;
wire \top/processor/sha_core/n3517_143 ;
wire \top/processor/sha_core/n3889_111 ;
wire \top/processor/sha_core/n3517_145 ;
wire \top/processor/sha_core/n3889_113 ;
wire \top/processor/sha_core/n3517_147 ;
wire \top/processor/sha_core/n3889_115 ;
wire \top/processor/sha_core/n3490_147 ;
wire \top/processor/sha_core/n3862_115 ;
wire \top/processor/sha_core/n3518_133 ;
wire \top/processor/sha_core/n3890_101 ;
wire \top/processor/sha_core/n3518_135 ;
wire \top/processor/sha_core/n3890_103 ;
wire \top/processor/sha_core/n3518_137 ;
wire \top/processor/sha_core/n3890_105 ;
wire \top/processor/sha_core/n3518_139 ;
wire \top/processor/sha_core/n3890_107 ;
wire \top/processor/sha_core/n3518_141 ;
wire \top/processor/sha_core/n3890_109 ;
wire \top/processor/sha_core/n3518_143 ;
wire \top/processor/sha_core/n3890_111 ;
wire \top/processor/sha_core/n3518_145 ;
wire \top/processor/sha_core/n3890_113 ;
wire \top/processor/sha_core/n3518_147 ;
wire \top/processor/sha_core/n3890_115 ;
wire \top/processor/sha_core/n3519_133 ;
wire \top/processor/sha_core/n3891_101 ;
wire \top/processor/sha_core/n3519_135 ;
wire \top/processor/sha_core/n3891_103 ;
wire \top/processor/sha_core/n3491_133 ;
wire \top/processor/sha_core/n3863_101 ;
wire \top/processor/sha_core/n3519_137 ;
wire \top/processor/sha_core/n3891_105 ;
wire \top/processor/sha_core/n3519_139 ;
wire \top/processor/sha_core/n3891_107 ;
wire \top/processor/sha_core/n3519_141 ;
wire \top/processor/sha_core/n3891_109 ;
wire \top/processor/sha_core/n3519_143 ;
wire \top/processor/sha_core/n3891_111 ;
wire \top/processor/sha_core/n3519_145 ;
wire \top/processor/sha_core/n3891_113 ;
wire \top/processor/sha_core/n3519_147 ;
wire \top/processor/sha_core/n3891_115 ;
wire \top/processor/sha_core/n3607_149 ;
wire \top/processor/sha_core/n3608_149 ;
wire \top/processor/sha_core/n3609_149 ;
wire \top/processor/sha_core/n3610_149 ;
wire \top/processor/sha_core/n3611_149 ;
wire \top/processor/sha_core/n3612_149 ;
wire \top/processor/sha_core/n3613_149 ;
wire \top/processor/sha_core/n3491_135 ;
wire \top/processor/sha_core/n3863_103 ;
wire \top/processor/sha_core/n3614_149 ;
wire \top/processor/sha_core/n3615_149 ;
wire \top/processor/sha_core/n3616_149 ;
wire \top/processor/sha_core/n3617_149 ;
wire \top/processor/sha_core/n3618_149 ;
wire \top/processor/sha_core/n3619_149 ;
wire \top/processor/sha_core/n3620_149 ;
wire \top/processor/sha_core/n3621_149 ;
wire \top/processor/sha_core/n3622_149 ;
wire \top/processor/sha_core/n3623_149 ;
wire \top/processor/sha_core/n3624_149 ;
wire \top/processor/sha_core/n3625_149 ;
wire \top/processor/sha_core/n3626_149 ;
wire \top/processor/sha_core/n3627_149 ;
wire \top/processor/sha_core/n3628_149 ;
wire \top/processor/sha_core/n3629_149 ;
wire \top/processor/sha_core/n3630_149 ;
wire \top/processor/sha_core/n3631_149 ;
wire \top/processor/sha_core/n3632_149 ;
wire \top/processor/sha_core/n3633_149 ;
wire \top/processor/sha_core/n3491_137 ;
wire \top/processor/sha_core/n3863_105 ;
wire \top/processor/sha_core/n3634_149 ;
wire \top/processor/sha_core/n3635_149 ;
wire \top/processor/sha_core/n3636_149 ;
wire \top/processor/sha_core/n3637_149 ;
wire \top/processor/sha_core/n3638_149 ;
wire \top/processor/sha_core/n3491_139 ;
wire \top/processor/sha_core/n3863_107 ;
wire \top/processor/sha_core/n3607_151 ;
wire \top/processor/sha_core/n3608_151 ;
wire \top/processor/sha_core/n3609_151 ;
wire \top/processor/sha_core/n3491_141 ;
wire \top/processor/sha_core/n3863_109 ;
wire \top/processor/sha_core/n3610_151 ;
wire \top/processor/sha_core/n3611_151 ;
wire \top/processor/sha_core/n3612_151 ;
wire \top/processor/sha_core/n3613_151 ;
wire \top/processor/sha_core/n3614_151 ;
wire \top/processor/sha_core/n3615_151 ;
wire \top/processor/sha_core/n3616_151 ;
wire \top/processor/sha_core/n3617_151 ;
wire \top/processor/sha_core/n3618_151 ;
wire \top/processor/sha_core/n3619_151 ;
wire \top/processor/sha_core/n3620_151 ;
wire \top/processor/sha_core/n3621_151 ;
wire \top/processor/sha_core/n3622_151 ;
wire \top/processor/sha_core/n3623_151 ;
wire \top/processor/sha_core/n3624_151 ;
wire \top/processor/sha_core/n3625_151 ;
wire \top/processor/sha_core/n3626_151 ;
wire \top/processor/sha_core/n3627_151 ;
wire \top/processor/sha_core/n3628_151 ;
wire \top/processor/sha_core/n3629_151 ;
wire \top/processor/sha_core/n3491_143 ;
wire \top/processor/sha_core/n3863_111 ;
wire \top/processor/sha_core/n3488_143 ;
wire \top/processor/sha_core/n3860_111 ;
wire \top/processor/sha_core/n3630_151 ;
wire \top/processor/sha_core/n3631_151 ;
wire \top/processor/sha_core/n3632_151 ;
wire \top/processor/sha_core/n3633_151 ;
wire \top/processor/sha_core/n3634_151 ;
wire \top/processor/sha_core/n3635_151 ;
wire \top/processor/sha_core/n3636_151 ;
wire \top/processor/sha_core/n3637_151 ;
wire \top/processor/sha_core/n3638_151 ;
wire \top/processor/sha_core/n3491_145 ;
wire \top/processor/sha_core/n3863_113 ;
wire \top/processor/sha_core/n3491_147 ;
wire \top/processor/sha_core/n3863_115 ;
wire \top/processor/sha_core/n3607_153 ;
wire \top/processor/sha_core/n3608_153 ;
wire \top/processor/sha_core/n3609_153 ;
wire \top/processor/sha_core/n3610_153 ;
wire \top/processor/sha_core/n3611_153 ;
wire \top/processor/sha_core/n3612_153 ;
wire \top/processor/sha_core/n3613_153 ;
wire \top/processor/sha_core/n3614_153 ;
wire \top/processor/sha_core/n3615_153 ;
wire \top/processor/sha_core/n3616_153 ;
wire \top/processor/sha_core/n3617_153 ;
wire \top/processor/sha_core/n3618_153 ;
wire \top/processor/sha_core/n3619_153 ;
wire \top/processor/sha_core/n3620_153 ;
wire \top/processor/sha_core/n3621_153 ;
wire \top/processor/sha_core/n3622_153 ;
wire \top/processor/sha_core/n3623_153 ;
wire \top/processor/sha_core/n3624_153 ;
wire \top/processor/sha_core/n3625_153 ;
wire \top/processor/sha_core/n3492_133 ;
wire \top/processor/sha_core/n3864_101 ;
wire \top/processor/sha_core/n3626_153 ;
wire \top/processor/sha_core/n3627_153 ;
wire \top/processor/sha_core/n3628_153 ;
wire \top/processor/sha_core/n3629_153 ;
wire \top/processor/sha_core/n3630_153 ;
wire \top/processor/sha_core/n3631_153 ;
wire \top/processor/sha_core/n3632_153 ;
wire \top/processor/sha_core/n3633_153 ;
wire \top/processor/sha_core/n3634_153 ;
wire \top/processor/sha_core/n3635_153 ;
wire \top/processor/sha_core/n3636_153 ;
wire \top/processor/sha_core/n3637_153 ;
wire \top/processor/sha_core/n3638_153 ;
wire \top/processor/sha_core/n3492_135 ;
wire \top/processor/sha_core/n3864_103 ;
wire \top/processor/sha_core/n3492_137 ;
wire \top/processor/sha_core/n3864_105 ;
wire \top/processor/sha_core/n3607_155 ;
wire \top/processor/sha_core/n3608_155 ;
wire \top/processor/sha_core/n3609_155 ;
wire \top/processor/sha_core/n3610_155 ;
wire \top/processor/sha_core/n3611_155 ;
wire \top/processor/sha_core/n3612_155 ;
wire \top/processor/sha_core/n3613_155 ;
wire \top/processor/sha_core/n3614_155 ;
wire \top/processor/sha_core/n3615_155 ;
wire \top/processor/sha_core/n3616_155 ;
wire \top/processor/sha_core/n3617_155 ;
wire \top/processor/sha_core/n3618_155 ;
wire \top/processor/sha_core/n3619_155 ;
wire \top/processor/sha_core/n3620_155 ;
wire \top/processor/sha_core/n3621_155 ;
wire \top/processor/sha_core/n3492_139 ;
wire \top/processor/sha_core/n3864_107 ;
wire \top/processor/sha_core/n3622_155 ;
wire \top/processor/sha_core/n3623_155 ;
wire \top/processor/sha_core/n3624_155 ;
wire \top/processor/sha_core/n3625_155 ;
wire \top/processor/sha_core/n3626_155 ;
wire \top/processor/sha_core/n3627_155 ;
wire \top/processor/sha_core/n3628_155 ;
wire \top/processor/sha_core/n3629_155 ;
wire \top/processor/sha_core/n3630_155 ;
wire \top/processor/sha_core/n3631_155 ;
wire \top/processor/sha_core/n3632_155 ;
wire \top/processor/sha_core/n3633_155 ;
wire \top/processor/sha_core/n3634_155 ;
wire \top/processor/sha_core/n3635_155 ;
wire \top/processor/sha_core/n3636_155 ;
wire \top/processor/sha_core/n3637_155 ;
wire \top/processor/sha_core/n3638_155 ;
wire \top/processor/sha_core/n3492_141 ;
wire \top/processor/sha_core/n3864_109 ;
wire \top/processor/sha_core/n3492_143 ;
wire \top/processor/sha_core/n3864_111 ;
wire \top/processor/sha_core/n3607_157 ;
wire \top/processor/sha_core/n3608_157 ;
wire \top/processor/sha_core/n3609_157 ;
wire \top/processor/sha_core/n3610_157 ;
wire \top/processor/sha_core/n3611_157 ;
wire \top/processor/sha_core/n3612_157 ;
wire \top/processor/sha_core/n3613_157 ;
wire \top/processor/sha_core/n3614_157 ;
wire \top/processor/sha_core/n3615_157 ;
wire \top/processor/sha_core/n3616_157 ;
wire \top/processor/sha_core/n3617_157 ;
wire \top/processor/sha_core/n3492_145 ;
wire \top/processor/sha_core/n3864_113 ;
wire \top/processor/sha_core/n3618_157 ;
wire \top/processor/sha_core/n3619_157 ;
wire \top/processor/sha_core/n3620_157 ;
wire \top/processor/sha_core/n3621_157 ;
wire \top/processor/sha_core/n3622_157 ;
wire \top/processor/sha_core/n3623_157 ;
wire \top/processor/sha_core/n3624_157 ;
wire \top/processor/sha_core/n3625_157 ;
wire \top/processor/sha_core/n3626_157 ;
wire \top/processor/sha_core/n3627_157 ;
wire \top/processor/sha_core/n3628_157 ;
wire \top/processor/sha_core/n3629_157 ;
wire \top/processor/sha_core/n3630_157 ;
wire \top/processor/sha_core/n3631_157 ;
wire \top/processor/sha_core/n3632_157 ;
wire \top/processor/sha_core/n3633_157 ;
wire \top/processor/sha_core/n3634_157 ;
wire \top/processor/sha_core/n3635_157 ;
wire \top/processor/sha_core/n3636_157 ;
wire \top/processor/sha_core/n3637_157 ;
wire \top/processor/sha_core/n3492_147 ;
wire \top/processor/sha_core/n3864_115 ;
wire \top/processor/sha_core/n3488_145 ;
wire \top/processor/sha_core/n3860_113 ;
wire \top/processor/sha_core/n3638_157 ;
wire \top/processor/sha_core/n3493_133 ;
wire \top/processor/sha_core/n3865_101 ;
wire \top/processor/sha_core/n3607_159 ;
wire \top/processor/sha_core/n3608_159 ;
wire \top/processor/sha_core/n3609_159 ;
wire \top/processor/sha_core/n3610_159 ;
wire \top/processor/sha_core/n3611_159 ;
wire \top/processor/sha_core/n3612_159 ;
wire \top/processor/sha_core/n3613_159 ;
wire \top/processor/sha_core/n3493_135 ;
wire \top/processor/sha_core/n3865_103 ;
wire \top/processor/sha_core/n3614_159 ;
wire \top/processor/sha_core/n3615_159 ;
wire \top/processor/sha_core/n3616_159 ;
wire \top/processor/sha_core/n3617_159 ;
wire \top/processor/sha_core/n3618_159 ;
wire \top/processor/sha_core/n3619_159 ;
wire \top/processor/sha_core/n3620_159 ;
wire \top/processor/sha_core/n3621_159 ;
wire \top/processor/sha_core/n3622_159 ;
wire \top/processor/sha_core/n3623_159 ;
wire \top/processor/sha_core/n3624_159 ;
wire \top/processor/sha_core/n3625_159 ;
wire \top/processor/sha_core/n3626_159 ;
wire \top/processor/sha_core/n3627_159 ;
wire \top/processor/sha_core/n3628_159 ;
wire \top/processor/sha_core/n3629_159 ;
wire \top/processor/sha_core/n3630_159 ;
wire \top/processor/sha_core/n3631_159 ;
wire \top/processor/sha_core/n3632_159 ;
wire \top/processor/sha_core/n3633_159 ;
wire \top/processor/sha_core/n3493_137 ;
wire \top/processor/sha_core/n3865_105 ;
wire \top/processor/sha_core/n3634_159 ;
wire \top/processor/sha_core/n3635_159 ;
wire \top/processor/sha_core/n3636_159 ;
wire \top/processor/sha_core/n3637_159 ;
wire \top/processor/sha_core/n3638_159 ;
wire \top/processor/sha_core/n3493_139 ;
wire \top/processor/sha_core/n3865_107 ;
wire \top/processor/sha_core/n3607_161 ;
wire \top/processor/sha_core/n3608_161 ;
wire \top/processor/sha_core/n3609_161 ;
wire \top/processor/sha_core/n3493_141 ;
wire \top/processor/sha_core/n3865_109 ;
wire \top/processor/sha_core/n3610_161 ;
wire \top/processor/sha_core/n3611_161 ;
wire \top/processor/sha_core/n3612_161 ;
wire \top/processor/sha_core/n3613_161 ;
wire \top/processor/sha_core/n3614_161 ;
wire \top/processor/sha_core/n3615_161 ;
wire \top/processor/sha_core/n3616_161 ;
wire \top/processor/sha_core/n3617_161 ;
wire \top/processor/sha_core/n3618_161 ;
wire \top/processor/sha_core/n3619_161 ;
wire \top/processor/sha_core/n3620_161 ;
wire \top/processor/sha_core/n3621_161 ;
wire \top/processor/sha_core/n3622_161 ;
wire \top/processor/sha_core/n3623_161 ;
wire \top/processor/sha_core/n3624_161 ;
wire \top/processor/sha_core/n3625_161 ;
wire \top/processor/sha_core/n3626_161 ;
wire \top/processor/sha_core/n3627_161 ;
wire \top/processor/sha_core/n3628_161 ;
wire \top/processor/sha_core/n3629_161 ;
wire \top/processor/sha_core/n3493_143 ;
wire \top/processor/sha_core/n3865_111 ;
wire \top/processor/sha_core/n3630_161 ;
wire \top/processor/sha_core/n3631_161 ;
wire \top/processor/sha_core/n3632_161 ;
wire \top/processor/sha_core/n3633_161 ;
wire \top/processor/sha_core/n3634_161 ;
wire \top/processor/sha_core/n3635_161 ;
wire \top/processor/sha_core/n3636_161 ;
wire \top/processor/sha_core/n3637_161 ;
wire \top/processor/sha_core/n3638_161 ;
wire \top/processor/sha_core/n3493_145 ;
wire \top/processor/sha_core/n3865_113 ;
wire \top/processor/sha_core/n3493_147 ;
wire \top/processor/sha_core/n3865_115 ;
wire \top/processor/sha_core/n3607_163 ;
wire \top/processor/sha_core/n3608_163 ;
wire \top/processor/sha_core/n3609_163 ;
wire \top/processor/sha_core/n3610_163 ;
wire \top/processor/sha_core/n3611_163 ;
wire \top/processor/sha_core/n3612_163 ;
wire \top/processor/sha_core/n3613_163 ;
wire \top/processor/sha_core/n3614_163 ;
wire \top/processor/sha_core/n3615_163 ;
wire \top/processor/sha_core/n3616_163 ;
wire \top/processor/sha_core/n3617_163 ;
wire \top/processor/sha_core/n3618_163 ;
wire \top/processor/sha_core/n3619_163 ;
wire \top/processor/sha_core/n3620_163 ;
wire \top/processor/sha_core/n3621_163 ;
wire \top/processor/sha_core/n3622_163 ;
wire \top/processor/sha_core/n3623_163 ;
wire \top/processor/sha_core/n3624_163 ;
wire \top/processor/sha_core/n3625_163 ;
wire \top/processor/sha_core/n3494_145 ;
wire \top/processor/sha_core/n3866_113 ;
wire \top/processor/sha_core/n3626_163 ;
wire \top/processor/sha_core/n3627_163 ;
wire \top/processor/sha_core/n3628_163 ;
wire \top/processor/sha_core/n3629_163 ;
wire \top/processor/sha_core/n3630_163 ;
wire \top/processor/sha_core/n3631_163 ;
wire \top/processor/sha_core/n3632_163 ;
wire \top/processor/sha_core/n3633_163 ;
wire \top/processor/sha_core/n3634_163 ;
wire \top/processor/sha_core/n3635_163 ;
wire \top/processor/sha_core/n3636_163 ;
wire \top/processor/sha_core/n3637_163 ;
wire \top/processor/sha_core/n3638_163 ;
wire \top/processor/sha_core/n3494_147 ;
wire \top/processor/sha_core/n3866_115 ;
wire \top/processor/sha_core/n3488_147 ;
wire \top/processor/sha_core/n3860_115 ;
wire \top/processor/sha_core/n3494_149 ;
wire \top/processor/sha_core/n3494_150 ;
wire \top/processor/sha_core/n3494_151 ;
wire \top/processor/sha_core/n3866_116 ;
wire \top/processor/sha_core/n3866_117 ;
wire \top/processor/sha_core/n3607_164 ;
wire \top/processor/sha_core/n3608_164 ;
wire \top/processor/sha_core/n3609_164 ;
wire \top/processor/sha_core/n3610_164 ;
wire \top/processor/sha_core/n3611_164 ;
wire \top/processor/sha_core/n3612_164 ;
wire \top/processor/sha_core/n3613_164 ;
wire \top/processor/sha_core/n3614_164 ;
wire \top/processor/sha_core/n3615_164 ;
wire \top/processor/sha_core/n3616_164 ;
wire \top/processor/sha_core/n3617_164 ;
wire \top/processor/sha_core/n3618_164 ;
wire \top/processor/sha_core/n3619_164 ;
wire \top/processor/sha_core/n3620_164 ;
wire \top/processor/sha_core/n3621_164 ;
wire \top/processor/sha_core/n3494_152 ;
wire \top/processor/sha_core/n3494_153 ;
wire \top/processor/sha_core/n3494_154 ;
wire \top/processor/sha_core/n3866_118 ;
wire \top/processor/sha_core/n3866_119 ;
wire \top/processor/sha_core/n3622_164 ;
wire \top/processor/sha_core/n3623_164 ;
wire \top/processor/sha_core/n3624_164 ;
wire \top/processor/sha_core/n3625_164 ;
wire \top/processor/sha_core/n3626_164 ;
wire \top/processor/sha_core/n3627_164 ;
wire \top/processor/sha_core/n3628_164 ;
wire \top/processor/sha_core/n3629_164 ;
wire \top/processor/sha_core/n3630_164 ;
wire \top/processor/sha_core/n3631_164 ;
wire \top/processor/sha_core/n3632_164 ;
wire \top/processor/sha_core/n3633_164 ;
wire \top/processor/sha_core/n3634_164 ;
wire \top/processor/sha_core/n3635_164 ;
wire \top/processor/sha_core/n3636_164 ;
wire \top/processor/sha_core/n3637_164 ;
wire \top/processor/sha_core/n3638_164 ;
wire \top/processor/sha_core/n3494_155 ;
wire \top/processor/sha_core/n3494_156 ;
wire \top/processor/sha_core/n3494_157 ;
wire \top/processor/sha_core/n3866_120 ;
wire \top/processor/sha_core/n3866_121 ;
wire \top/processor/sha_core/n3494_158 ;
wire \top/processor/sha_core/n3494_159 ;
wire \top/processor/sha_core/n3494_160 ;
wire \top/processor/sha_core/n3866_122 ;
wire \top/processor/sha_core/n3866_123 ;
wire \top/processor/sha_core/n3607_165 ;
wire \top/processor/sha_core/n3608_165 ;
wire \top/processor/sha_core/n3609_165 ;
wire \top/processor/sha_core/n3610_165 ;
wire \top/processor/sha_core/n3611_165 ;
wire \top/processor/sha_core/n3612_165 ;
wire \top/processor/sha_core/n3613_165 ;
wire \top/processor/sha_core/n3614_165 ;
wire \top/processor/sha_core/n3615_165 ;
wire \top/processor/sha_core/n3616_165 ;
wire \top/processor/sha_core/n3617_165 ;
wire \top/processor/sha_core/n3494_161 ;
wire \top/processor/sha_core/n3494_162 ;
wire \top/processor/sha_core/n3494_163 ;
wire \top/processor/sha_core/n3866_124 ;
wire \top/processor/sha_core/n3866_125 ;
wire \top/processor/sha_core/n3618_165 ;
wire \top/processor/sha_core/n3619_165 ;
wire \top/processor/sha_core/n3620_165 ;
wire \top/processor/sha_core/n3621_165 ;
wire \top/processor/sha_core/n3622_165 ;
wire \top/processor/sha_core/n3623_165 ;
wire \top/processor/sha_core/n3624_165 ;
wire \top/processor/sha_core/n3625_165 ;
wire \top/processor/sha_core/n3626_165 ;
wire \top/processor/sha_core/n3627_165 ;
wire \top/processor/sha_core/n3628_165 ;
wire \top/processor/sha_core/n3629_165 ;
wire \top/processor/sha_core/n3630_165 ;
wire \top/processor/sha_core/n3631_165 ;
wire \top/processor/sha_core/n3632_165 ;
wire \top/processor/sha_core/n3633_165 ;
wire \top/processor/sha_core/n3634_165 ;
wire \top/processor/sha_core/n3635_165 ;
wire \top/processor/sha_core/n3636_165 ;
wire \top/processor/sha_core/n3637_165 ;
wire \top/processor/sha_core/n3494_164 ;
wire \top/processor/sha_core/n3494_165 ;
wire \top/processor/sha_core/n3494_166 ;
wire \top/processor/sha_core/n3866_126 ;
wire \top/processor/sha_core/n3866_127 ;
wire \top/processor/sha_core/n3638_165 ;
wire \top/processor/sha_core/n3495_148 ;
wire \top/processor/sha_core/n3495_149 ;
wire \top/processor/sha_core/n3495_150 ;
wire \top/processor/sha_core/n3867_116 ;
wire \top/processor/sha_core/n3867_117 ;
wire \top/processor/sha_core/n3607_166 ;
wire \top/processor/sha_core/n3608_166 ;
wire \top/processor/sha_core/n3609_166 ;
wire \top/processor/sha_core/n3610_166 ;
wire \top/processor/sha_core/n3611_166 ;
wire \top/processor/sha_core/n3612_166 ;
wire \top/processor/sha_core/n3613_166 ;
wire \top/processor/sha_core/n3495_151 ;
wire \top/processor/sha_core/n3495_152 ;
wire \top/processor/sha_core/n3495_153 ;
wire \top/processor/sha_core/n3867_118 ;
wire \top/processor/sha_core/n3867_119 ;
wire \top/processor/sha_core/n3614_166 ;
wire \top/processor/sha_core/n3615_166 ;
wire \top/processor/sha_core/n3616_166 ;
wire \top/processor/sha_core/n3617_166 ;
wire \top/processor/sha_core/n3618_166 ;
wire \top/processor/sha_core/n3619_166 ;
wire \top/processor/sha_core/n3620_166 ;
wire \top/processor/sha_core/n3621_166 ;
wire \top/processor/sha_core/n3622_166 ;
wire \top/processor/sha_core/n3623_166 ;
wire \top/processor/sha_core/n3624_166 ;
wire \top/processor/sha_core/n3625_166 ;
wire \top/processor/sha_core/n3626_166 ;
wire \top/processor/sha_core/n3627_166 ;
wire \top/processor/sha_core/n3628_166 ;
wire \top/processor/sha_core/n3629_166 ;
wire \top/processor/sha_core/n3630_166 ;
wire \top/processor/sha_core/n3631_166 ;
wire \top/processor/sha_core/n3632_166 ;
wire \top/processor/sha_core/n3633_166 ;
wire \top/processor/sha_core/n3495_154 ;
wire \top/processor/sha_core/n3495_155 ;
wire \top/processor/sha_core/n3495_156 ;
wire \top/processor/sha_core/n3867_120 ;
wire \top/processor/sha_core/n3867_121 ;
wire \top/processor/sha_core/n3634_166 ;
wire \top/processor/sha_core/n3635_166 ;
wire \top/processor/sha_core/n3636_166 ;
wire \top/processor/sha_core/n3637_166 ;
wire \top/processor/sha_core/n3638_166 ;
wire \top/processor/sha_core/n3495_157 ;
wire \top/processor/sha_core/n3495_158 ;
wire \top/processor/sha_core/n3495_159 ;
wire \top/processor/sha_core/n3867_122 ;
wire \top/processor/sha_core/n3867_123 ;
wire \top/processor/sha_core/n3488_148 ;
wire \top/processor/sha_core/n3488_149 ;
wire \top/processor/sha_core/n3488_150 ;
wire \top/processor/sha_core/n3860_116 ;
wire \top/processor/sha_core/n3860_117 ;
wire \top/processor/sha_core/n3607_167 ;
wire \top/processor/sha_core/n3608_167 ;
wire \top/processor/sha_core/n3609_167 ;
wire \top/processor/sha_core/n3495_160 ;
wire \top/processor/sha_core/n3495_161 ;
wire \top/processor/sha_core/n3495_162 ;
wire \top/processor/sha_core/n3867_124 ;
wire \top/processor/sha_core/n3867_125 ;
wire \top/processor/sha_core/n3610_167 ;
wire \top/processor/sha_core/n3611_167 ;
wire \top/processor/sha_core/n3612_167 ;
wire \top/processor/sha_core/n3613_167 ;
wire \top/processor/sha_core/n3614_167 ;
wire \top/processor/sha_core/n3615_167 ;
wire \top/processor/sha_core/n3616_167 ;
wire \top/processor/sha_core/n3617_167 ;
wire \top/processor/sha_core/n3618_167 ;
wire \top/processor/sha_core/n3619_167 ;
wire \top/processor/sha_core/n3620_167 ;
wire \top/processor/sha_core/n3621_167 ;
wire \top/processor/sha_core/n3622_167 ;
wire \top/processor/sha_core/n3623_167 ;
wire \top/processor/sha_core/n3624_167 ;
wire \top/processor/sha_core/n3625_167 ;
wire \top/processor/sha_core/n3626_167 ;
wire \top/processor/sha_core/n3627_167 ;
wire \top/processor/sha_core/n3628_167 ;
wire \top/processor/sha_core/n3629_167 ;
wire \top/processor/sha_core/n3495_163 ;
wire \top/processor/sha_core/n3495_164 ;
wire \top/processor/sha_core/n3495_165 ;
wire \top/processor/sha_core/n3867_126 ;
wire \top/processor/sha_core/n3867_127 ;
wire \top/processor/sha_core/n3630_167 ;
wire \top/processor/sha_core/n3631_167 ;
wire \top/processor/sha_core/n3632_167 ;
wire \top/processor/sha_core/n3633_167 ;
wire \top/processor/sha_core/n3634_167 ;
wire \top/processor/sha_core/n3635_167 ;
wire \top/processor/sha_core/n3636_167 ;
wire \top/processor/sha_core/n3637_167 ;
wire \top/processor/sha_core/n3638_167 ;
wire \top/processor/sha_core/n3495_166 ;
wire \top/processor/sha_core/n3495_167 ;
wire \top/processor/sha_core/n3495_168 ;
wire \top/processor/sha_core/n3867_128 ;
wire \top/processor/sha_core/n3867_129 ;
wire \top/processor/sha_core/n3495_169 ;
wire \top/processor/sha_core/n3495_170 ;
wire \top/processor/sha_core/n3495_171 ;
wire \top/processor/sha_core/n3867_130 ;
wire \top/processor/sha_core/n3867_131 ;
wire \top/processor/sha_core/n3607_168 ;
wire \top/processor/sha_core/n3608_168 ;
wire \top/processor/sha_core/n3609_168 ;
wire \top/processor/sha_core/n3610_168 ;
wire \top/processor/sha_core/n3611_168 ;
wire \top/processor/sha_core/n3612_168 ;
wire \top/processor/sha_core/n3613_168 ;
wire \top/processor/sha_core/n3614_168 ;
wire \top/processor/sha_core/n3615_168 ;
wire \top/processor/sha_core/n3616_168 ;
wire \top/processor/sha_core/n3617_168 ;
wire \top/processor/sha_core/n3618_168 ;
wire \top/processor/sha_core/n3619_168 ;
wire \top/processor/sha_core/n3620_168 ;
wire \top/processor/sha_core/n3621_168 ;
wire \top/processor/sha_core/n3622_168 ;
wire \top/processor/sha_core/n3623_168 ;
wire \top/processor/sha_core/n3624_168 ;
wire \top/processor/sha_core/n3625_168 ;
wire \top/processor/sha_core/n3496_148 ;
wire \top/processor/sha_core/n3496_149 ;
wire \top/processor/sha_core/n3496_150 ;
wire \top/processor/sha_core/n3868_116 ;
wire \top/processor/sha_core/n3868_117 ;
wire \top/processor/sha_core/n3626_168 ;
wire \top/processor/sha_core/n3627_168 ;
wire \top/processor/sha_core/n3628_168 ;
wire \top/processor/sha_core/n3629_168 ;
wire \top/processor/sha_core/n3630_168 ;
wire \top/processor/sha_core/n3631_168 ;
wire \top/processor/sha_core/n3632_168 ;
wire \top/processor/sha_core/n3633_168 ;
wire \top/processor/sha_core/n3634_168 ;
wire \top/processor/sha_core/n3635_168 ;
wire \top/processor/sha_core/n3636_168 ;
wire \top/processor/sha_core/n3637_168 ;
wire \top/processor/sha_core/n3638_168 ;
wire \top/processor/sha_core/n3496_151 ;
wire \top/processor/sha_core/n3496_152 ;
wire \top/processor/sha_core/n3496_153 ;
wire \top/processor/sha_core/n3868_118 ;
wire \top/processor/sha_core/n3868_119 ;
wire \top/processor/sha_core/n3496_154 ;
wire \top/processor/sha_core/n3496_155 ;
wire \top/processor/sha_core/n3496_156 ;
wire \top/processor/sha_core/n3868_120 ;
wire \top/processor/sha_core/n3868_121 ;
wire \top/processor/sha_core/n3607_169 ;
wire \top/processor/sha_core/n3608_169 ;
wire \top/processor/sha_core/n3609_169 ;
wire \top/processor/sha_core/n3610_169 ;
wire \top/processor/sha_core/n3611_169 ;
wire \top/processor/sha_core/n3612_169 ;
wire \top/processor/sha_core/n3613_169 ;
wire \top/processor/sha_core/n3614_169 ;
wire \top/processor/sha_core/n3615_169 ;
wire \top/processor/sha_core/n3616_169 ;
wire \top/processor/sha_core/n3617_169 ;
wire \top/processor/sha_core/n3618_169 ;
wire \top/processor/sha_core/n3619_169 ;
wire \top/processor/sha_core/n3620_169 ;
wire \top/processor/sha_core/n3621_169 ;
wire \top/processor/sha_core/n3496_157 ;
wire \top/processor/sha_core/n3496_158 ;
wire \top/processor/sha_core/n3496_159 ;
wire \top/processor/sha_core/n3868_122 ;
wire \top/processor/sha_core/n3868_123 ;
wire \top/processor/sha_core/n3622_169 ;
wire \top/processor/sha_core/n3623_169 ;
wire \top/processor/sha_core/n3624_169 ;
wire \top/processor/sha_core/n3625_169 ;
wire \top/processor/sha_core/n3626_169 ;
wire \top/processor/sha_core/n3627_169 ;
wire \top/processor/sha_core/n3628_169 ;
wire \top/processor/sha_core/n3629_169 ;
wire \top/processor/sha_core/n3630_169 ;
wire \top/processor/sha_core/n3631_169 ;
wire \top/processor/sha_core/n3632_169 ;
wire \top/processor/sha_core/n3633_169 ;
wire \top/processor/sha_core/n3634_169 ;
wire \top/processor/sha_core/n3635_169 ;
wire \top/processor/sha_core/n3636_169 ;
wire \top/processor/sha_core/n3637_169 ;
wire \top/processor/sha_core/n3638_169 ;
wire \top/processor/sha_core/n3496_160 ;
wire \top/processor/sha_core/n3496_161 ;
wire \top/processor/sha_core/n3496_162 ;
wire \top/processor/sha_core/n3868_124 ;
wire \top/processor/sha_core/n3868_125 ;
wire \top/processor/sha_core/n3496_163 ;
wire \top/processor/sha_core/n3496_164 ;
wire \top/processor/sha_core/n3496_165 ;
wire \top/processor/sha_core/n3868_126 ;
wire \top/processor/sha_core/n3868_127 ;
wire \top/processor/sha_core/n3488_151 ;
wire \top/processor/sha_core/n3488_152 ;
wire \top/processor/sha_core/n3488_153 ;
wire \top/processor/sha_core/n3860_118 ;
wire \top/processor/sha_core/n3860_119 ;
wire \top/processor/sha_core/n3607_170 ;
wire \top/processor/sha_core/n3608_170 ;
wire \top/processor/sha_core/n3609_170 ;
wire \top/processor/sha_core/n3610_170 ;
wire \top/processor/sha_core/n3611_170 ;
wire \top/processor/sha_core/n3612_170 ;
wire \top/processor/sha_core/n3613_170 ;
wire \top/processor/sha_core/n3614_170 ;
wire \top/processor/sha_core/n3615_170 ;
wire \top/processor/sha_core/n3616_170 ;
wire \top/processor/sha_core/n3617_170 ;
wire \top/processor/sha_core/n3496_166 ;
wire \top/processor/sha_core/n3496_167 ;
wire \top/processor/sha_core/n3496_168 ;
wire \top/processor/sha_core/n3868_128 ;
wire \top/processor/sha_core/n3868_129 ;
wire \top/processor/sha_core/n3618_170 ;
wire \top/processor/sha_core/n3619_170 ;
wire \top/processor/sha_core/n3620_170 ;
wire \top/processor/sha_core/n3621_170 ;
wire \top/processor/sha_core/n3622_170 ;
wire \top/processor/sha_core/n3623_170 ;
wire \top/processor/sha_core/n3624_170 ;
wire \top/processor/sha_core/n3625_170 ;
wire \top/processor/sha_core/n3626_170 ;
wire \top/processor/sha_core/n3627_170 ;
wire \top/processor/sha_core/n3628_170 ;
wire \top/processor/sha_core/n3629_170 ;
wire \top/processor/sha_core/n3630_170 ;
wire \top/processor/sha_core/n3631_170 ;
wire \top/processor/sha_core/n3632_170 ;
wire \top/processor/sha_core/n3633_170 ;
wire \top/processor/sha_core/n3634_170 ;
wire \top/processor/sha_core/n3635_170 ;
wire \top/processor/sha_core/n3636_170 ;
wire \top/processor/sha_core/n3637_170 ;
wire \top/processor/sha_core/n3496_169 ;
wire \top/processor/sha_core/n3496_170 ;
wire \top/processor/sha_core/n3496_171 ;
wire \top/processor/sha_core/n3868_130 ;
wire \top/processor/sha_core/n3868_131 ;
wire \top/processor/sha_core/n3638_170 ;
wire \top/processor/sha_core/n3497_148 ;
wire \top/processor/sha_core/n3497_149 ;
wire \top/processor/sha_core/n3497_150 ;
wire \top/processor/sha_core/n3869_116 ;
wire \top/processor/sha_core/n3869_117 ;
wire \top/processor/sha_core/n3607_171 ;
wire \top/processor/sha_core/n3608_171 ;
wire \top/processor/sha_core/n3609_171 ;
wire \top/processor/sha_core/n3610_171 ;
wire \top/processor/sha_core/n3611_171 ;
wire \top/processor/sha_core/n3612_171 ;
wire \top/processor/sha_core/n3613_171 ;
wire \top/processor/sha_core/n3497_151 ;
wire \top/processor/sha_core/n3497_152 ;
wire \top/processor/sha_core/n3497_153 ;
wire \top/processor/sha_core/n3869_118 ;
wire \top/processor/sha_core/n3869_119 ;
wire \top/processor/sha_core/n3614_171 ;
wire \top/processor/sha_core/n3615_171 ;
wire \top/processor/sha_core/n3616_171 ;
wire \top/processor/sha_core/n3617_171 ;
wire \top/processor/sha_core/n3618_171 ;
wire \top/processor/sha_core/n3619_171 ;
wire \top/processor/sha_core/n3620_171 ;
wire \top/processor/sha_core/n3621_171 ;
wire \top/processor/sha_core/n3622_171 ;
wire \top/processor/sha_core/n3623_171 ;
wire \top/processor/sha_core/n3624_171 ;
wire \top/processor/sha_core/n3625_171 ;
wire \top/processor/sha_core/n3626_171 ;
wire \top/processor/sha_core/n3627_171 ;
wire \top/processor/sha_core/n3628_171 ;
wire \top/processor/sha_core/n3629_171 ;
wire \top/processor/sha_core/n3630_171 ;
wire \top/processor/sha_core/n3631_171 ;
wire \top/processor/sha_core/n3632_171 ;
wire \top/processor/sha_core/n3633_171 ;
wire \top/processor/sha_core/n3497_154 ;
wire \top/processor/sha_core/n3497_155 ;
wire \top/processor/sha_core/n3497_156 ;
wire \top/processor/sha_core/n3869_120 ;
wire \top/processor/sha_core/n3869_121 ;
wire \top/processor/sha_core/n3634_171 ;
wire \top/processor/sha_core/n3635_171 ;
wire \top/processor/sha_core/n3636_171 ;
wire \top/processor/sha_core/n3637_171 ;
wire \top/processor/sha_core/n3638_171 ;
wire \top/processor/sha_core/n3497_157 ;
wire \top/processor/sha_core/n3497_158 ;
wire \top/processor/sha_core/n3497_159 ;
wire \top/processor/sha_core/n3869_122 ;
wire \top/processor/sha_core/n3869_123 ;
wire \top/processor/sha_core/n3497_160 ;
wire \top/processor/sha_core/n3497_161 ;
wire \top/processor/sha_core/n3497_162 ;
wire \top/processor/sha_core/n3869_124 ;
wire \top/processor/sha_core/n3869_125 ;
wire \top/processor/sha_core/n3497_163 ;
wire \top/processor/sha_core/n3497_164 ;
wire \top/processor/sha_core/n3497_165 ;
wire \top/processor/sha_core/n3869_126 ;
wire \top/processor/sha_core/n3869_127 ;
wire \top/processor/sha_core/n3497_166 ;
wire \top/processor/sha_core/n3497_167 ;
wire \top/processor/sha_core/n3497_168 ;
wire \top/processor/sha_core/n3869_128 ;
wire \top/processor/sha_core/n3869_129 ;
wire \top/processor/sha_core/n3497_169 ;
wire \top/processor/sha_core/n3497_170 ;
wire \top/processor/sha_core/n3497_171 ;
wire \top/processor/sha_core/n3869_130 ;
wire \top/processor/sha_core/n3869_131 ;
wire \top/processor/sha_core/n3488_154 ;
wire \top/processor/sha_core/n3488_155 ;
wire \top/processor/sha_core/n3488_156 ;
wire \top/processor/sha_core/n3860_120 ;
wire \top/processor/sha_core/n3860_121 ;
wire \top/processor/sha_core/n3498_148 ;
wire \top/processor/sha_core/n3498_149 ;
wire \top/processor/sha_core/n3498_150 ;
wire \top/processor/sha_core/n3870_116 ;
wire \top/processor/sha_core/n3870_117 ;
wire \top/processor/sha_core/n3498_151 ;
wire \top/processor/sha_core/n3498_152 ;
wire \top/processor/sha_core/n3498_153 ;
wire \top/processor/sha_core/n3870_118 ;
wire \top/processor/sha_core/n3870_119 ;
wire \top/processor/sha_core/n3498_154 ;
wire \top/processor/sha_core/n3498_155 ;
wire \top/processor/sha_core/n3498_156 ;
wire \top/processor/sha_core/n3870_120 ;
wire \top/processor/sha_core/n3870_121 ;
wire \top/processor/sha_core/n3498_157 ;
wire \top/processor/sha_core/n3498_158 ;
wire \top/processor/sha_core/n3498_159 ;
wire \top/processor/sha_core/n3870_122 ;
wire \top/processor/sha_core/n3870_123 ;
wire \top/processor/sha_core/n3498_160 ;
wire \top/processor/sha_core/n3498_161 ;
wire \top/processor/sha_core/n3498_162 ;
wire \top/processor/sha_core/n3870_124 ;
wire \top/processor/sha_core/n3870_125 ;
wire \top/processor/sha_core/n3498_163 ;
wire \top/processor/sha_core/n3498_164 ;
wire \top/processor/sha_core/n3498_165 ;
wire \top/processor/sha_core/n3870_126 ;
wire \top/processor/sha_core/n3870_127 ;
wire \top/processor/sha_core/n3498_166 ;
wire \top/processor/sha_core/n3498_167 ;
wire \top/processor/sha_core/n3498_168 ;
wire \top/processor/sha_core/n3870_128 ;
wire \top/processor/sha_core/n3870_129 ;
wire \top/processor/sha_core/n3498_169 ;
wire \top/processor/sha_core/n3498_170 ;
wire \top/processor/sha_core/n3498_171 ;
wire \top/processor/sha_core/n3870_130 ;
wire \top/processor/sha_core/n3870_131 ;
wire \top/processor/sha_core/n3499_148 ;
wire \top/processor/sha_core/n3499_149 ;
wire \top/processor/sha_core/n3499_150 ;
wire \top/processor/sha_core/n3871_116 ;
wire \top/processor/sha_core/n3871_117 ;
wire \top/processor/sha_core/n3499_151 ;
wire \top/processor/sha_core/n3499_152 ;
wire \top/processor/sha_core/n3499_153 ;
wire \top/processor/sha_core/n3871_118 ;
wire \top/processor/sha_core/n3871_119 ;
wire \top/processor/sha_core/n3489_148 ;
wire \top/processor/sha_core/n3489_149 ;
wire \top/processor/sha_core/n3489_150 ;
wire \top/processor/sha_core/n3861_116 ;
wire \top/processor/sha_core/n3861_117 ;
wire \top/processor/sha_core/n3499_154 ;
wire \top/processor/sha_core/n3499_155 ;
wire \top/processor/sha_core/n3499_156 ;
wire \top/processor/sha_core/n3871_120 ;
wire \top/processor/sha_core/n3871_121 ;
wire \top/processor/sha_core/n3499_157 ;
wire \top/processor/sha_core/n3499_158 ;
wire \top/processor/sha_core/n3499_159 ;
wire \top/processor/sha_core/n3871_122 ;
wire \top/processor/sha_core/n3871_123 ;
wire \top/processor/sha_core/n3499_160 ;
wire \top/processor/sha_core/n3499_161 ;
wire \top/processor/sha_core/n3499_162 ;
wire \top/processor/sha_core/n3871_124 ;
wire \top/processor/sha_core/n3871_125 ;
wire \top/processor/sha_core/n3499_163 ;
wire \top/processor/sha_core/n3499_164 ;
wire \top/processor/sha_core/n3499_165 ;
wire \top/processor/sha_core/n3871_126 ;
wire \top/processor/sha_core/n3871_127 ;
wire \top/processor/sha_core/n3499_166 ;
wire \top/processor/sha_core/n3499_167 ;
wire \top/processor/sha_core/n3499_168 ;
wire \top/processor/sha_core/n3871_128 ;
wire \top/processor/sha_core/n3871_129 ;
wire \top/processor/sha_core/n3499_169 ;
wire \top/processor/sha_core/n3499_170 ;
wire \top/processor/sha_core/n3499_171 ;
wire \top/processor/sha_core/n3871_130 ;
wire \top/processor/sha_core/n3871_131 ;
wire \top/processor/sha_core/n3500_148 ;
wire \top/processor/sha_core/n3500_149 ;
wire \top/processor/sha_core/n3500_150 ;
wire \top/processor/sha_core/n3872_116 ;
wire \top/processor/sha_core/n3872_117 ;
wire \top/processor/sha_core/n3500_151 ;
wire \top/processor/sha_core/n3500_152 ;
wire \top/processor/sha_core/n3500_153 ;
wire \top/processor/sha_core/n3872_118 ;
wire \top/processor/sha_core/n3872_119 ;
wire \top/processor/sha_core/n3500_154 ;
wire \top/processor/sha_core/n3500_155 ;
wire \top/processor/sha_core/n3500_156 ;
wire \top/processor/sha_core/n3872_120 ;
wire \top/processor/sha_core/n3872_121 ;
wire \top/processor/sha_core/n3500_157 ;
wire \top/processor/sha_core/n3500_158 ;
wire \top/processor/sha_core/n3500_159 ;
wire \top/processor/sha_core/n3872_122 ;
wire \top/processor/sha_core/n3872_123 ;
wire \top/processor/sha_core/n3489_151 ;
wire \top/processor/sha_core/n3489_152 ;
wire \top/processor/sha_core/n3489_153 ;
wire \top/processor/sha_core/n3861_118 ;
wire \top/processor/sha_core/n3861_119 ;
wire \top/processor/sha_core/n3488_157 ;
wire \top/processor/sha_core/n3488_158 ;
wire \top/processor/sha_core/n3488_159 ;
wire \top/processor/sha_core/n3860_122 ;
wire \top/processor/sha_core/n3860_123 ;
wire \top/processor/sha_core/n3500_160 ;
wire \top/processor/sha_core/n3500_161 ;
wire \top/processor/sha_core/n3500_162 ;
wire \top/processor/sha_core/n3872_124 ;
wire \top/processor/sha_core/n3872_125 ;
wire \top/processor/sha_core/n3500_163 ;
wire \top/processor/sha_core/n3500_164 ;
wire \top/processor/sha_core/n3500_165 ;
wire \top/processor/sha_core/n3872_126 ;
wire \top/processor/sha_core/n3872_127 ;
wire \top/processor/sha_core/n3500_166 ;
wire \top/processor/sha_core/n3500_167 ;
wire \top/processor/sha_core/n3500_168 ;
wire \top/processor/sha_core/n3872_128 ;
wire \top/processor/sha_core/n3872_129 ;
wire \top/processor/sha_core/n3500_169 ;
wire \top/processor/sha_core/n3500_170 ;
wire \top/processor/sha_core/n3500_171 ;
wire \top/processor/sha_core/n3872_130 ;
wire \top/processor/sha_core/n3872_131 ;
wire \top/processor/sha_core/n3501_148 ;
wire \top/processor/sha_core/n3501_149 ;
wire \top/processor/sha_core/n3501_150 ;
wire \top/processor/sha_core/n3873_116 ;
wire \top/processor/sha_core/n3873_117 ;
wire \top/processor/sha_core/n3501_151 ;
wire \top/processor/sha_core/n3501_152 ;
wire \top/processor/sha_core/n3501_153 ;
wire \top/processor/sha_core/n3873_118 ;
wire \top/processor/sha_core/n3873_119 ;
wire \top/processor/sha_core/n3501_154 ;
wire \top/processor/sha_core/n3501_155 ;
wire \top/processor/sha_core/n3501_156 ;
wire \top/processor/sha_core/n3873_120 ;
wire \top/processor/sha_core/n3873_121 ;
wire \top/processor/sha_core/n3501_157 ;
wire \top/processor/sha_core/n3501_158 ;
wire \top/processor/sha_core/n3501_159 ;
wire \top/processor/sha_core/n3873_122 ;
wire \top/processor/sha_core/n3873_123 ;
wire \top/processor/sha_core/n3501_160 ;
wire \top/processor/sha_core/n3501_161 ;
wire \top/processor/sha_core/n3501_162 ;
wire \top/processor/sha_core/n3873_124 ;
wire \top/processor/sha_core/n3873_125 ;
wire \top/processor/sha_core/n3501_163 ;
wire \top/processor/sha_core/n3501_164 ;
wire \top/processor/sha_core/n3501_165 ;
wire \top/processor/sha_core/n3873_126 ;
wire \top/processor/sha_core/n3873_127 ;
wire \top/processor/sha_core/n3489_154 ;
wire \top/processor/sha_core/n3489_155 ;
wire \top/processor/sha_core/n3489_156 ;
wire \top/processor/sha_core/n3861_120 ;
wire \top/processor/sha_core/n3861_121 ;
wire \top/processor/sha_core/n3501_166 ;
wire \top/processor/sha_core/n3501_167 ;
wire \top/processor/sha_core/n3501_168 ;
wire \top/processor/sha_core/n3873_128 ;
wire \top/processor/sha_core/n3873_129 ;
wire \top/processor/sha_core/n3501_169 ;
wire \top/processor/sha_core/n3501_170 ;
wire \top/processor/sha_core/n3501_171 ;
wire \top/processor/sha_core/n3873_130 ;
wire \top/processor/sha_core/n3873_131 ;
wire \top/processor/sha_core/n3502_148 ;
wire \top/processor/sha_core/n3502_149 ;
wire \top/processor/sha_core/n3502_150 ;
wire \top/processor/sha_core/n3874_116 ;
wire \top/processor/sha_core/n3874_117 ;
wire \top/processor/sha_core/n3502_151 ;
wire \top/processor/sha_core/n3502_152 ;
wire \top/processor/sha_core/n3502_153 ;
wire \top/processor/sha_core/n3874_118 ;
wire \top/processor/sha_core/n3874_119 ;
wire \top/processor/sha_core/n3502_154 ;
wire \top/processor/sha_core/n3502_155 ;
wire \top/processor/sha_core/n3502_156 ;
wire \top/processor/sha_core/n3874_120 ;
wire \top/processor/sha_core/n3874_121 ;
wire \top/processor/sha_core/n3502_157 ;
wire \top/processor/sha_core/n3502_158 ;
wire \top/processor/sha_core/n3502_159 ;
wire \top/processor/sha_core/n3874_122 ;
wire \top/processor/sha_core/n3874_123 ;
wire \top/processor/sha_core/n3502_160 ;
wire \top/processor/sha_core/n3502_161 ;
wire \top/processor/sha_core/n3502_162 ;
wire \top/processor/sha_core/n3874_124 ;
wire \top/processor/sha_core/n3874_125 ;
wire \top/processor/sha_core/n3502_163 ;
wire \top/processor/sha_core/n3502_164 ;
wire \top/processor/sha_core/n3502_165 ;
wire \top/processor/sha_core/n3874_126 ;
wire \top/processor/sha_core/n3874_127 ;
wire \top/processor/sha_core/n3502_166 ;
wire \top/processor/sha_core/n3502_167 ;
wire \top/processor/sha_core/n3502_168 ;
wire \top/processor/sha_core/n3874_128 ;
wire \top/processor/sha_core/n3874_129 ;
wire \top/processor/sha_core/n3502_169 ;
wire \top/processor/sha_core/n3502_170 ;
wire \top/processor/sha_core/n3502_171 ;
wire \top/processor/sha_core/n3874_130 ;
wire \top/processor/sha_core/n3874_131 ;
wire \top/processor/sha_core/n3489_157 ;
wire \top/processor/sha_core/n3489_158 ;
wire \top/processor/sha_core/n3489_159 ;
wire \top/processor/sha_core/n3861_122 ;
wire \top/processor/sha_core/n3861_123 ;
wire \top/processor/sha_core/n3503_148 ;
wire \top/processor/sha_core/n3503_149 ;
wire \top/processor/sha_core/n3503_150 ;
wire \top/processor/sha_core/n3875_116 ;
wire \top/processor/sha_core/n3875_117 ;
wire \top/processor/sha_core/n3503_151 ;
wire \top/processor/sha_core/n3503_152 ;
wire \top/processor/sha_core/n3503_153 ;
wire \top/processor/sha_core/n3875_118 ;
wire \top/processor/sha_core/n3875_119 ;
wire \top/processor/sha_core/n3503_154 ;
wire \top/processor/sha_core/n3503_155 ;
wire \top/processor/sha_core/n3503_156 ;
wire \top/processor/sha_core/n3875_120 ;
wire \top/processor/sha_core/n3875_121 ;
wire \top/processor/sha_core/n3503_157 ;
wire \top/processor/sha_core/n3503_158 ;
wire \top/processor/sha_core/n3503_159 ;
wire \top/processor/sha_core/n3875_122 ;
wire \top/processor/sha_core/n3875_123 ;
wire \top/processor/sha_core/n3503_160 ;
wire \top/processor/sha_core/n3503_161 ;
wire \top/processor/sha_core/n3503_162 ;
wire \top/processor/sha_core/n3875_124 ;
wire \top/processor/sha_core/n3875_125 ;
wire \top/processor/sha_core/n3503_163 ;
wire \top/processor/sha_core/n3503_164 ;
wire \top/processor/sha_core/n3503_165 ;
wire \top/processor/sha_core/n3875_126 ;
wire \top/processor/sha_core/n3875_127 ;
wire \top/processor/sha_core/n3503_166 ;
wire \top/processor/sha_core/n3503_167 ;
wire \top/processor/sha_core/n3503_168 ;
wire \top/processor/sha_core/n3875_128 ;
wire \top/processor/sha_core/n3875_129 ;
wire \top/processor/sha_core/n3503_169 ;
wire \top/processor/sha_core/n3503_170 ;
wire \top/processor/sha_core/n3503_171 ;
wire \top/processor/sha_core/n3875_130 ;
wire \top/processor/sha_core/n3875_131 ;
wire \top/processor/sha_core/n3504_148 ;
wire \top/processor/sha_core/n3504_149 ;
wire \top/processor/sha_core/n3504_150 ;
wire \top/processor/sha_core/n3876_116 ;
wire \top/processor/sha_core/n3876_117 ;
wire \top/processor/sha_core/n3504_151 ;
wire \top/processor/sha_core/n3504_152 ;
wire \top/processor/sha_core/n3504_153 ;
wire \top/processor/sha_core/n3876_118 ;
wire \top/processor/sha_core/n3876_119 ;
wire \top/processor/sha_core/n3489_160 ;
wire \top/processor/sha_core/n3489_161 ;
wire \top/processor/sha_core/n3489_162 ;
wire \top/processor/sha_core/n3861_124 ;
wire \top/processor/sha_core/n3861_125 ;
wire \top/processor/sha_core/n3504_154 ;
wire \top/processor/sha_core/n3504_155 ;
wire \top/processor/sha_core/n3504_156 ;
wire \top/processor/sha_core/n3876_120 ;
wire \top/processor/sha_core/n3876_121 ;
wire \top/processor/sha_core/n3504_157 ;
wire \top/processor/sha_core/n3504_158 ;
wire \top/processor/sha_core/n3504_159 ;
wire \top/processor/sha_core/n3876_122 ;
wire \top/processor/sha_core/n3876_123 ;
wire \top/processor/sha_core/n3504_160 ;
wire \top/processor/sha_core/n3504_161 ;
wire \top/processor/sha_core/n3504_162 ;
wire \top/processor/sha_core/n3876_124 ;
wire \top/processor/sha_core/n3876_125 ;
wire \top/processor/sha_core/n3504_163 ;
wire \top/processor/sha_core/n3504_164 ;
wire \top/processor/sha_core/n3504_165 ;
wire \top/processor/sha_core/n3876_126 ;
wire \top/processor/sha_core/n3876_127 ;
wire \top/processor/sha_core/n3504_166 ;
wire \top/processor/sha_core/n3504_167 ;
wire \top/processor/sha_core/n3504_168 ;
wire \top/processor/sha_core/n3876_128 ;
wire \top/processor/sha_core/n3876_129 ;
wire \top/processor/sha_core/n3504_169 ;
wire \top/processor/sha_core/n3504_170 ;
wire \top/processor/sha_core/n3504_171 ;
wire \top/processor/sha_core/n3876_130 ;
wire \top/processor/sha_core/n3876_131 ;
wire \top/processor/sha_core/n3505_148 ;
wire \top/processor/sha_core/n3505_149 ;
wire \top/processor/sha_core/n3505_150 ;
wire \top/processor/sha_core/n3877_116 ;
wire \top/processor/sha_core/n3877_117 ;
wire \top/processor/sha_core/n3505_151 ;
wire \top/processor/sha_core/n3505_152 ;
wire \top/processor/sha_core/n3505_153 ;
wire \top/processor/sha_core/n3877_118 ;
wire \top/processor/sha_core/n3877_119 ;
wire \top/processor/sha_core/n3505_154 ;
wire \top/processor/sha_core/n3505_155 ;
wire \top/processor/sha_core/n3505_156 ;
wire \top/processor/sha_core/n3877_120 ;
wire \top/processor/sha_core/n3877_121 ;
wire \top/processor/sha_core/n3505_157 ;
wire \top/processor/sha_core/n3505_158 ;
wire \top/processor/sha_core/n3505_159 ;
wire \top/processor/sha_core/n3877_122 ;
wire \top/processor/sha_core/n3877_123 ;
wire \top/processor/sha_core/n3489_163 ;
wire \top/processor/sha_core/n3489_164 ;
wire \top/processor/sha_core/n3489_165 ;
wire \top/processor/sha_core/n3861_126 ;
wire \top/processor/sha_core/n3861_127 ;
wire \top/processor/sha_core/n3505_160 ;
wire \top/processor/sha_core/n3505_161 ;
wire \top/processor/sha_core/n3505_162 ;
wire \top/processor/sha_core/n3877_124 ;
wire \top/processor/sha_core/n3877_125 ;
wire \top/processor/sha_core/n3505_163 ;
wire \top/processor/sha_core/n3505_164 ;
wire \top/processor/sha_core/n3505_165 ;
wire \top/processor/sha_core/n3877_126 ;
wire \top/processor/sha_core/n3877_127 ;
wire \top/processor/sha_core/n3505_166 ;
wire \top/processor/sha_core/n3505_167 ;
wire \top/processor/sha_core/n3505_168 ;
wire \top/processor/sha_core/n3877_128 ;
wire \top/processor/sha_core/n3877_129 ;
wire \top/processor/sha_core/n3505_169 ;
wire \top/processor/sha_core/n3505_170 ;
wire \top/processor/sha_core/n3505_171 ;
wire \top/processor/sha_core/n3877_130 ;
wire \top/processor/sha_core/n3877_131 ;
wire \top/processor/sha_core/n3506_148 ;
wire \top/processor/sha_core/n3506_149 ;
wire \top/processor/sha_core/n3506_150 ;
wire \top/processor/sha_core/n3878_116 ;
wire \top/processor/sha_core/n3878_117 ;
wire \top/processor/sha_core/n3506_151 ;
wire \top/processor/sha_core/n3506_152 ;
wire \top/processor/sha_core/n3506_153 ;
wire \top/processor/sha_core/n3878_118 ;
wire \top/processor/sha_core/n3878_119 ;
wire \top/processor/sha_core/n3506_154 ;
wire \top/processor/sha_core/n3506_155 ;
wire \top/processor/sha_core/n3506_156 ;
wire \top/processor/sha_core/n3878_120 ;
wire \top/processor/sha_core/n3878_121 ;
wire \top/processor/sha_core/n3506_157 ;
wire \top/processor/sha_core/n3506_158 ;
wire \top/processor/sha_core/n3506_159 ;
wire \top/processor/sha_core/n3878_122 ;
wire \top/processor/sha_core/n3878_123 ;
wire \top/processor/sha_core/n3506_160 ;
wire \top/processor/sha_core/n3506_161 ;
wire \top/processor/sha_core/n3506_162 ;
wire \top/processor/sha_core/n3878_124 ;
wire \top/processor/sha_core/n3878_125 ;
wire \top/processor/sha_core/n3506_163 ;
wire \top/processor/sha_core/n3506_164 ;
wire \top/processor/sha_core/n3506_165 ;
wire \top/processor/sha_core/n3878_126 ;
wire \top/processor/sha_core/n3878_127 ;
wire \top/processor/sha_core/n3489_166 ;
wire \top/processor/sha_core/n3489_167 ;
wire \top/processor/sha_core/n3489_168 ;
wire \top/processor/sha_core/n3861_128 ;
wire \top/processor/sha_core/n3861_129 ;
wire \top/processor/sha_core/n3506_166 ;
wire \top/processor/sha_core/n3506_167 ;
wire \top/processor/sha_core/n3506_168 ;
wire \top/processor/sha_core/n3878_128 ;
wire \top/processor/sha_core/n3878_129 ;
wire \top/processor/sha_core/n3506_169 ;
wire \top/processor/sha_core/n3506_170 ;
wire \top/processor/sha_core/n3506_171 ;
wire \top/processor/sha_core/n3878_130 ;
wire \top/processor/sha_core/n3878_131 ;
wire \top/processor/sha_core/n3507_148 ;
wire \top/processor/sha_core/n3507_149 ;
wire \top/processor/sha_core/n3507_150 ;
wire \top/processor/sha_core/n3879_116 ;
wire \top/processor/sha_core/n3879_117 ;
wire \top/processor/sha_core/n3507_151 ;
wire \top/processor/sha_core/n3507_152 ;
wire \top/processor/sha_core/n3507_153 ;
wire \top/processor/sha_core/n3879_118 ;
wire \top/processor/sha_core/n3879_119 ;
wire \top/processor/sha_core/n3507_154 ;
wire \top/processor/sha_core/n3507_155 ;
wire \top/processor/sha_core/n3507_156 ;
wire \top/processor/sha_core/n3879_120 ;
wire \top/processor/sha_core/n3879_121 ;
wire \top/processor/sha_core/n3507_157 ;
wire \top/processor/sha_core/n3507_158 ;
wire \top/processor/sha_core/n3507_159 ;
wire \top/processor/sha_core/n3879_122 ;
wire \top/processor/sha_core/n3879_123 ;
wire \top/processor/sha_core/n3507_160 ;
wire \top/processor/sha_core/n3507_161 ;
wire \top/processor/sha_core/n3507_162 ;
wire \top/processor/sha_core/n3879_124 ;
wire \top/processor/sha_core/n3879_125 ;
wire \top/processor/sha_core/n3507_163 ;
wire \top/processor/sha_core/n3507_164 ;
wire \top/processor/sha_core/n3507_165 ;
wire \top/processor/sha_core/n3879_126 ;
wire \top/processor/sha_core/n3879_127 ;
wire \top/processor/sha_core/n3507_166 ;
wire \top/processor/sha_core/n3507_167 ;
wire \top/processor/sha_core/n3507_168 ;
wire \top/processor/sha_core/n3879_128 ;
wire \top/processor/sha_core/n3879_129 ;
wire \top/processor/sha_core/n3507_169 ;
wire \top/processor/sha_core/n3507_170 ;
wire \top/processor/sha_core/n3507_171 ;
wire \top/processor/sha_core/n3879_130 ;
wire \top/processor/sha_core/n3879_131 ;
wire \top/processor/sha_core/n3489_169 ;
wire \top/processor/sha_core/n3489_170 ;
wire \top/processor/sha_core/n3489_171 ;
wire \top/processor/sha_core/n3861_130 ;
wire \top/processor/sha_core/n3861_131 ;
wire \top/processor/sha_core/n3508_148 ;
wire \top/processor/sha_core/n3508_149 ;
wire \top/processor/sha_core/n3508_150 ;
wire \top/processor/sha_core/n3880_116 ;
wire \top/processor/sha_core/n3880_117 ;
wire \top/processor/sha_core/n3508_151 ;
wire \top/processor/sha_core/n3508_152 ;
wire \top/processor/sha_core/n3508_153 ;
wire \top/processor/sha_core/n3880_118 ;
wire \top/processor/sha_core/n3880_119 ;
wire \top/processor/sha_core/n3508_154 ;
wire \top/processor/sha_core/n3508_155 ;
wire \top/processor/sha_core/n3508_156 ;
wire \top/processor/sha_core/n3880_120 ;
wire \top/processor/sha_core/n3880_121 ;
wire \top/processor/sha_core/n3508_157 ;
wire \top/processor/sha_core/n3508_158 ;
wire \top/processor/sha_core/n3508_159 ;
wire \top/processor/sha_core/n3880_122 ;
wire \top/processor/sha_core/n3880_123 ;
wire \top/processor/sha_core/n3508_160 ;
wire \top/processor/sha_core/n3508_161 ;
wire \top/processor/sha_core/n3508_162 ;
wire \top/processor/sha_core/n3880_124 ;
wire \top/processor/sha_core/n3880_125 ;
wire \top/processor/sha_core/n3508_163 ;
wire \top/processor/sha_core/n3508_164 ;
wire \top/processor/sha_core/n3508_165 ;
wire \top/processor/sha_core/n3880_126 ;
wire \top/processor/sha_core/n3880_127 ;
wire \top/processor/sha_core/n3508_166 ;
wire \top/processor/sha_core/n3508_167 ;
wire \top/processor/sha_core/n3508_168 ;
wire \top/processor/sha_core/n3880_128 ;
wire \top/processor/sha_core/n3880_129 ;
wire \top/processor/sha_core/n3508_169 ;
wire \top/processor/sha_core/n3508_170 ;
wire \top/processor/sha_core/n3508_171 ;
wire \top/processor/sha_core/n3880_130 ;
wire \top/processor/sha_core/n3880_131 ;
wire \top/processor/sha_core/n3509_148 ;
wire \top/processor/sha_core/n3509_149 ;
wire \top/processor/sha_core/n3509_150 ;
wire \top/processor/sha_core/n3881_116 ;
wire \top/processor/sha_core/n3881_117 ;
wire \top/processor/sha_core/n3509_151 ;
wire \top/processor/sha_core/n3509_152 ;
wire \top/processor/sha_core/n3509_153 ;
wire \top/processor/sha_core/n3881_118 ;
wire \top/processor/sha_core/n3881_119 ;
wire \top/processor/sha_core/n3490_148 ;
wire \top/processor/sha_core/n3490_149 ;
wire \top/processor/sha_core/n3490_150 ;
wire \top/processor/sha_core/n3862_116 ;
wire \top/processor/sha_core/n3862_117 ;
wire \top/processor/sha_core/n3509_154 ;
wire \top/processor/sha_core/n3509_155 ;
wire \top/processor/sha_core/n3509_156 ;
wire \top/processor/sha_core/n3881_120 ;
wire \top/processor/sha_core/n3881_121 ;
wire \top/processor/sha_core/n3509_157 ;
wire \top/processor/sha_core/n3509_158 ;
wire \top/processor/sha_core/n3509_159 ;
wire \top/processor/sha_core/n3881_122 ;
wire \top/processor/sha_core/n3881_123 ;
wire \top/processor/sha_core/n3509_160 ;
wire \top/processor/sha_core/n3509_161 ;
wire \top/processor/sha_core/n3509_162 ;
wire \top/processor/sha_core/n3881_124 ;
wire \top/processor/sha_core/n3881_125 ;
wire \top/processor/sha_core/n3509_163 ;
wire \top/processor/sha_core/n3509_164 ;
wire \top/processor/sha_core/n3509_165 ;
wire \top/processor/sha_core/n3881_126 ;
wire \top/processor/sha_core/n3881_127 ;
wire \top/processor/sha_core/n3509_166 ;
wire \top/processor/sha_core/n3509_167 ;
wire \top/processor/sha_core/n3509_168 ;
wire \top/processor/sha_core/n3881_128 ;
wire \top/processor/sha_core/n3881_129 ;
wire \top/processor/sha_core/n3509_169 ;
wire \top/processor/sha_core/n3509_170 ;
wire \top/processor/sha_core/n3509_171 ;
wire \top/processor/sha_core/n3881_130 ;
wire \top/processor/sha_core/n3881_131 ;
wire \top/processor/sha_core/n3510_148 ;
wire \top/processor/sha_core/n3510_149 ;
wire \top/processor/sha_core/n3510_150 ;
wire \top/processor/sha_core/n3882_116 ;
wire \top/processor/sha_core/n3882_117 ;
wire \top/processor/sha_core/n3510_151 ;
wire \top/processor/sha_core/n3510_152 ;
wire \top/processor/sha_core/n3510_153 ;
wire \top/processor/sha_core/n3882_118 ;
wire \top/processor/sha_core/n3882_119 ;
wire \top/processor/sha_core/n3510_154 ;
wire \top/processor/sha_core/n3510_155 ;
wire \top/processor/sha_core/n3510_156 ;
wire \top/processor/sha_core/n3882_120 ;
wire \top/processor/sha_core/n3882_121 ;
wire \top/processor/sha_core/n3510_157 ;
wire \top/processor/sha_core/n3510_158 ;
wire \top/processor/sha_core/n3510_159 ;
wire \top/processor/sha_core/n3882_122 ;
wire \top/processor/sha_core/n3882_123 ;
wire \top/processor/sha_core/n3490_151 ;
wire \top/processor/sha_core/n3490_152 ;
wire \top/processor/sha_core/n3490_153 ;
wire \top/processor/sha_core/n3862_118 ;
wire \top/processor/sha_core/n3862_119 ;
wire \top/processor/sha_core/n3510_160 ;
wire \top/processor/sha_core/n3510_161 ;
wire \top/processor/sha_core/n3510_162 ;
wire \top/processor/sha_core/n3882_124 ;
wire \top/processor/sha_core/n3882_125 ;
wire \top/processor/sha_core/n3510_163 ;
wire \top/processor/sha_core/n3510_164 ;
wire \top/processor/sha_core/n3510_165 ;
wire \top/processor/sha_core/n3882_126 ;
wire \top/processor/sha_core/n3882_127 ;
wire \top/processor/sha_core/n3510_166 ;
wire \top/processor/sha_core/n3510_167 ;
wire \top/processor/sha_core/n3510_168 ;
wire \top/processor/sha_core/n3882_128 ;
wire \top/processor/sha_core/n3882_129 ;
wire \top/processor/sha_core/n3510_169 ;
wire \top/processor/sha_core/n3510_170 ;
wire \top/processor/sha_core/n3510_171 ;
wire \top/processor/sha_core/n3882_130 ;
wire \top/processor/sha_core/n3882_131 ;
wire \top/processor/sha_core/n3511_148 ;
wire \top/processor/sha_core/n3511_149 ;
wire \top/processor/sha_core/n3511_150 ;
wire \top/processor/sha_core/n3883_116 ;
wire \top/processor/sha_core/n3883_117 ;
wire \top/processor/sha_core/n3511_151 ;
wire \top/processor/sha_core/n3511_152 ;
wire \top/processor/sha_core/n3511_153 ;
wire \top/processor/sha_core/n3883_118 ;
wire \top/processor/sha_core/n3883_119 ;
wire \top/processor/sha_core/n3511_154 ;
wire \top/processor/sha_core/n3511_155 ;
wire \top/processor/sha_core/n3511_156 ;
wire \top/processor/sha_core/n3883_120 ;
wire \top/processor/sha_core/n3883_121 ;
wire \top/processor/sha_core/n3511_157 ;
wire \top/processor/sha_core/n3511_158 ;
wire \top/processor/sha_core/n3511_159 ;
wire \top/processor/sha_core/n3883_122 ;
wire \top/processor/sha_core/n3883_123 ;
wire \top/processor/sha_core/n3511_160 ;
wire \top/processor/sha_core/n3511_161 ;
wire \top/processor/sha_core/n3511_162 ;
wire \top/processor/sha_core/n3883_124 ;
wire \top/processor/sha_core/n3883_125 ;
wire \top/processor/sha_core/n3511_163 ;
wire \top/processor/sha_core/n3511_164 ;
wire \top/processor/sha_core/n3511_165 ;
wire \top/processor/sha_core/n3883_126 ;
wire \top/processor/sha_core/n3883_127 ;
wire \top/processor/sha_core/n3490_154 ;
wire \top/processor/sha_core/n3490_155 ;
wire \top/processor/sha_core/n3490_156 ;
wire \top/processor/sha_core/n3862_120 ;
wire \top/processor/sha_core/n3862_121 ;
wire \top/processor/sha_core/n3511_166 ;
wire \top/processor/sha_core/n3511_167 ;
wire \top/processor/sha_core/n3511_168 ;
wire \top/processor/sha_core/n3883_128 ;
wire \top/processor/sha_core/n3883_129 ;
wire \top/processor/sha_core/n3511_169 ;
wire \top/processor/sha_core/n3511_170 ;
wire \top/processor/sha_core/n3511_171 ;
wire \top/processor/sha_core/n3883_130 ;
wire \top/processor/sha_core/n3883_131 ;
wire \top/processor/sha_core/n3512_148 ;
wire \top/processor/sha_core/n3512_149 ;
wire \top/processor/sha_core/n3512_150 ;
wire \top/processor/sha_core/n3884_116 ;
wire \top/processor/sha_core/n3884_117 ;
wire \top/processor/sha_core/n3512_151 ;
wire \top/processor/sha_core/n3512_152 ;
wire \top/processor/sha_core/n3512_153 ;
wire \top/processor/sha_core/n3884_118 ;
wire \top/processor/sha_core/n3884_119 ;
wire \top/processor/sha_core/n3512_154 ;
wire \top/processor/sha_core/n3512_155 ;
wire \top/processor/sha_core/n3512_156 ;
wire \top/processor/sha_core/n3884_120 ;
wire \top/processor/sha_core/n3884_121 ;
wire \top/processor/sha_core/n3512_157 ;
wire \top/processor/sha_core/n3512_158 ;
wire \top/processor/sha_core/n3512_159 ;
wire \top/processor/sha_core/n3884_122 ;
wire \top/processor/sha_core/n3884_123 ;
wire \top/processor/sha_core/n3512_160 ;
wire \top/processor/sha_core/n3512_161 ;
wire \top/processor/sha_core/n3512_162 ;
wire \top/processor/sha_core/n3884_124 ;
wire \top/processor/sha_core/n3884_125 ;
wire \top/processor/sha_core/n3512_163 ;
wire \top/processor/sha_core/n3512_164 ;
wire \top/processor/sha_core/n3512_165 ;
wire \top/processor/sha_core/n3884_126 ;
wire \top/processor/sha_core/n3884_127 ;
wire \top/processor/sha_core/n3512_166 ;
wire \top/processor/sha_core/n3512_167 ;
wire \top/processor/sha_core/n3512_168 ;
wire \top/processor/sha_core/n3884_128 ;
wire \top/processor/sha_core/n3884_129 ;
wire \top/processor/sha_core/n3512_169 ;
wire \top/processor/sha_core/n3512_170 ;
wire \top/processor/sha_core/n3512_171 ;
wire \top/processor/sha_core/n3884_130 ;
wire \top/processor/sha_core/n3884_131 ;
wire \top/processor/sha_core/n3490_157 ;
wire \top/processor/sha_core/n3490_158 ;
wire \top/processor/sha_core/n3490_159 ;
wire \top/processor/sha_core/n3862_122 ;
wire \top/processor/sha_core/n3862_123 ;
wire \top/processor/sha_core/n3488_160 ;
wire \top/processor/sha_core/n3488_161 ;
wire \top/processor/sha_core/n3488_162 ;
wire \top/processor/sha_core/n3860_124 ;
wire \top/processor/sha_core/n3860_125 ;
wire \top/processor/sha_core/n3513_148 ;
wire \top/processor/sha_core/n3513_149 ;
wire \top/processor/sha_core/n3513_150 ;
wire \top/processor/sha_core/n3885_116 ;
wire \top/processor/sha_core/n3885_117 ;
wire \top/processor/sha_core/n3513_151 ;
wire \top/processor/sha_core/n3513_152 ;
wire \top/processor/sha_core/n3513_153 ;
wire \top/processor/sha_core/n3885_118 ;
wire \top/processor/sha_core/n3885_119 ;
wire \top/processor/sha_core/n3513_154 ;
wire \top/processor/sha_core/n3513_155 ;
wire \top/processor/sha_core/n3513_156 ;
wire \top/processor/sha_core/n3885_120 ;
wire \top/processor/sha_core/n3885_121 ;
wire \top/processor/sha_core/n3513_157 ;
wire \top/processor/sha_core/n3513_158 ;
wire \top/processor/sha_core/n3513_159 ;
wire \top/processor/sha_core/n3885_122 ;
wire \top/processor/sha_core/n3885_123 ;
wire \top/processor/sha_core/n3513_160 ;
wire \top/processor/sha_core/n3513_161 ;
wire \top/processor/sha_core/n3513_162 ;
wire \top/processor/sha_core/n3885_124 ;
wire \top/processor/sha_core/n3885_125 ;
wire \top/processor/sha_core/n3513_163 ;
wire \top/processor/sha_core/n3513_164 ;
wire \top/processor/sha_core/n3513_165 ;
wire \top/processor/sha_core/n3885_126 ;
wire \top/processor/sha_core/n3885_127 ;
wire \top/processor/sha_core/n3513_166 ;
wire \top/processor/sha_core/n3513_167 ;
wire \top/processor/sha_core/n3513_168 ;
wire \top/processor/sha_core/n3885_128 ;
wire \top/processor/sha_core/n3885_129 ;
wire \top/processor/sha_core/n3513_169 ;
wire \top/processor/sha_core/n3513_170 ;
wire \top/processor/sha_core/n3513_171 ;
wire \top/processor/sha_core/n3885_130 ;
wire \top/processor/sha_core/n3885_131 ;
wire \top/processor/sha_core/n3514_148 ;
wire \top/processor/sha_core/n3514_149 ;
wire \top/processor/sha_core/n3514_150 ;
wire \top/processor/sha_core/n3886_116 ;
wire \top/processor/sha_core/n3886_117 ;
wire \top/processor/sha_core/n3514_151 ;
wire \top/processor/sha_core/n3514_152 ;
wire \top/processor/sha_core/n3514_153 ;
wire \top/processor/sha_core/n3886_118 ;
wire \top/processor/sha_core/n3886_119 ;
wire \top/processor/sha_core/n3490_160 ;
wire \top/processor/sha_core/n3490_161 ;
wire \top/processor/sha_core/n3490_162 ;
wire \top/processor/sha_core/n3862_124 ;
wire \top/processor/sha_core/n3862_125 ;
wire \top/processor/sha_core/n3514_154 ;
wire \top/processor/sha_core/n3514_155 ;
wire \top/processor/sha_core/n3514_156 ;
wire \top/processor/sha_core/n3886_120 ;
wire \top/processor/sha_core/n3886_121 ;
wire \top/processor/sha_core/n3514_157 ;
wire \top/processor/sha_core/n3514_158 ;
wire \top/processor/sha_core/n3514_159 ;
wire \top/processor/sha_core/n3886_122 ;
wire \top/processor/sha_core/n3886_123 ;
wire \top/processor/sha_core/n3514_160 ;
wire \top/processor/sha_core/n3514_161 ;
wire \top/processor/sha_core/n3514_162 ;
wire \top/processor/sha_core/n3886_124 ;
wire \top/processor/sha_core/n3886_125 ;
wire \top/processor/sha_core/n3514_163 ;
wire \top/processor/sha_core/n3514_164 ;
wire \top/processor/sha_core/n3514_165 ;
wire \top/processor/sha_core/n3886_126 ;
wire \top/processor/sha_core/n3886_127 ;
wire \top/processor/sha_core/n3514_166 ;
wire \top/processor/sha_core/n3514_167 ;
wire \top/processor/sha_core/n3514_168 ;
wire \top/processor/sha_core/n3886_128 ;
wire \top/processor/sha_core/n3886_129 ;
wire \top/processor/sha_core/n3514_169 ;
wire \top/processor/sha_core/n3514_170 ;
wire \top/processor/sha_core/n3514_171 ;
wire \top/processor/sha_core/n3886_130 ;
wire \top/processor/sha_core/n3886_131 ;
wire \top/processor/sha_core/n3515_148 ;
wire \top/processor/sha_core/n3515_149 ;
wire \top/processor/sha_core/n3515_150 ;
wire \top/processor/sha_core/n3887_116 ;
wire \top/processor/sha_core/n3887_117 ;
wire \top/processor/sha_core/n3515_151 ;
wire \top/processor/sha_core/n3515_152 ;
wire \top/processor/sha_core/n3515_153 ;
wire \top/processor/sha_core/n3887_118 ;
wire \top/processor/sha_core/n3887_119 ;
wire \top/processor/sha_core/n3515_154 ;
wire \top/processor/sha_core/n3515_155 ;
wire \top/processor/sha_core/n3515_156 ;
wire \top/processor/sha_core/n3887_120 ;
wire \top/processor/sha_core/n3887_121 ;
wire \top/processor/sha_core/n3515_157 ;
wire \top/processor/sha_core/n3515_158 ;
wire \top/processor/sha_core/n3515_159 ;
wire \top/processor/sha_core/n3887_122 ;
wire \top/processor/sha_core/n3887_123 ;
wire \top/processor/sha_core/n3490_163 ;
wire \top/processor/sha_core/n3490_164 ;
wire \top/processor/sha_core/n3490_165 ;
wire \top/processor/sha_core/n3862_126 ;
wire \top/processor/sha_core/n3862_127 ;
wire \top/processor/sha_core/n3515_160 ;
wire \top/processor/sha_core/n3515_161 ;
wire \top/processor/sha_core/n3515_162 ;
wire \top/processor/sha_core/n3887_124 ;
wire \top/processor/sha_core/n3887_125 ;
wire \top/processor/sha_core/n3515_163 ;
wire \top/processor/sha_core/n3515_164 ;
wire \top/processor/sha_core/n3515_165 ;
wire \top/processor/sha_core/n3887_126 ;
wire \top/processor/sha_core/n3887_127 ;
wire \top/processor/sha_core/n3515_166 ;
wire \top/processor/sha_core/n3515_167 ;
wire \top/processor/sha_core/n3515_168 ;
wire \top/processor/sha_core/n3887_128 ;
wire \top/processor/sha_core/n3887_129 ;
wire \top/processor/sha_core/n3515_169 ;
wire \top/processor/sha_core/n3515_170 ;
wire \top/processor/sha_core/n3515_171 ;
wire \top/processor/sha_core/n3887_130 ;
wire \top/processor/sha_core/n3887_131 ;
wire \top/processor/sha_core/n3516_148 ;
wire \top/processor/sha_core/n3516_149 ;
wire \top/processor/sha_core/n3516_150 ;
wire \top/processor/sha_core/n3888_116 ;
wire \top/processor/sha_core/n3888_117 ;
wire \top/processor/sha_core/n3516_151 ;
wire \top/processor/sha_core/n3516_152 ;
wire \top/processor/sha_core/n3516_153 ;
wire \top/processor/sha_core/n3888_118 ;
wire \top/processor/sha_core/n3888_119 ;
wire \top/processor/sha_core/n3516_154 ;
wire \top/processor/sha_core/n3516_155 ;
wire \top/processor/sha_core/n3516_156 ;
wire \top/processor/sha_core/n3888_120 ;
wire \top/processor/sha_core/n3888_121 ;
wire \top/processor/sha_core/n3516_157 ;
wire \top/processor/sha_core/n3516_158 ;
wire \top/processor/sha_core/n3516_159 ;
wire \top/processor/sha_core/n3888_122 ;
wire \top/processor/sha_core/n3888_123 ;
wire \top/processor/sha_core/n3516_160 ;
wire \top/processor/sha_core/n3516_161 ;
wire \top/processor/sha_core/n3516_162 ;
wire \top/processor/sha_core/n3888_124 ;
wire \top/processor/sha_core/n3888_125 ;
wire \top/processor/sha_core/n3516_163 ;
wire \top/processor/sha_core/n3516_164 ;
wire \top/processor/sha_core/n3516_165 ;
wire \top/processor/sha_core/n3888_126 ;
wire \top/processor/sha_core/n3888_127 ;
wire \top/processor/sha_core/n3490_166 ;
wire \top/processor/sha_core/n3490_167 ;
wire \top/processor/sha_core/n3490_168 ;
wire \top/processor/sha_core/n3862_128 ;
wire \top/processor/sha_core/n3862_129 ;
wire \top/processor/sha_core/n3516_166 ;
wire \top/processor/sha_core/n3516_167 ;
wire \top/processor/sha_core/n3516_168 ;
wire \top/processor/sha_core/n3888_128 ;
wire \top/processor/sha_core/n3888_129 ;
wire \top/processor/sha_core/n3516_169 ;
wire \top/processor/sha_core/n3516_170 ;
wire \top/processor/sha_core/n3516_171 ;
wire \top/processor/sha_core/n3888_130 ;
wire \top/processor/sha_core/n3888_131 ;
wire \top/processor/sha_core/n3517_148 ;
wire \top/processor/sha_core/n3517_149 ;
wire \top/processor/sha_core/n3517_150 ;
wire \top/processor/sha_core/n3889_116 ;
wire \top/processor/sha_core/n3889_117 ;
wire \top/processor/sha_core/n3517_151 ;
wire \top/processor/sha_core/n3517_152 ;
wire \top/processor/sha_core/n3517_153 ;
wire \top/processor/sha_core/n3889_118 ;
wire \top/processor/sha_core/n3889_119 ;
wire \top/processor/sha_core/n3517_154 ;
wire \top/processor/sha_core/n3517_155 ;
wire \top/processor/sha_core/n3517_156 ;
wire \top/processor/sha_core/n3889_120 ;
wire \top/processor/sha_core/n3889_121 ;
wire \top/processor/sha_core/n3517_157 ;
wire \top/processor/sha_core/n3517_158 ;
wire \top/processor/sha_core/n3517_159 ;
wire \top/processor/sha_core/n3889_122 ;
wire \top/processor/sha_core/n3889_123 ;
wire \top/processor/sha_core/n3517_160 ;
wire \top/processor/sha_core/n3517_161 ;
wire \top/processor/sha_core/n3517_162 ;
wire \top/processor/sha_core/n3889_124 ;
wire \top/processor/sha_core/n3889_125 ;
wire \top/processor/sha_core/n3517_163 ;
wire \top/processor/sha_core/n3517_164 ;
wire \top/processor/sha_core/n3517_165 ;
wire \top/processor/sha_core/n3889_126 ;
wire \top/processor/sha_core/n3889_127 ;
wire \top/processor/sha_core/n3517_166 ;
wire \top/processor/sha_core/n3517_167 ;
wire \top/processor/sha_core/n3517_168 ;
wire \top/processor/sha_core/n3889_128 ;
wire \top/processor/sha_core/n3889_129 ;
wire \top/processor/sha_core/n3517_169 ;
wire \top/processor/sha_core/n3517_170 ;
wire \top/processor/sha_core/n3517_171 ;
wire \top/processor/sha_core/n3889_130 ;
wire \top/processor/sha_core/n3889_131 ;
wire \top/processor/sha_core/n3490_169 ;
wire \top/processor/sha_core/n3490_170 ;
wire \top/processor/sha_core/n3490_171 ;
wire \top/processor/sha_core/n3862_130 ;
wire \top/processor/sha_core/n3862_131 ;
wire \top/processor/sha_core/n3518_148 ;
wire \top/processor/sha_core/n3518_149 ;
wire \top/processor/sha_core/n3518_150 ;
wire \top/processor/sha_core/n3890_116 ;
wire \top/processor/sha_core/n3890_117 ;
wire \top/processor/sha_core/n3518_151 ;
wire \top/processor/sha_core/n3518_152 ;
wire \top/processor/sha_core/n3518_153 ;
wire \top/processor/sha_core/n3890_118 ;
wire \top/processor/sha_core/n3890_119 ;
wire \top/processor/sha_core/n3518_154 ;
wire \top/processor/sha_core/n3518_155 ;
wire \top/processor/sha_core/n3518_156 ;
wire \top/processor/sha_core/n3890_120 ;
wire \top/processor/sha_core/n3890_121 ;
wire \top/processor/sha_core/n3518_157 ;
wire \top/processor/sha_core/n3518_158 ;
wire \top/processor/sha_core/n3518_159 ;
wire \top/processor/sha_core/n3890_122 ;
wire \top/processor/sha_core/n3890_123 ;
wire \top/processor/sha_core/n3518_160 ;
wire \top/processor/sha_core/n3518_161 ;
wire \top/processor/sha_core/n3518_162 ;
wire \top/processor/sha_core/n3890_124 ;
wire \top/processor/sha_core/n3890_125 ;
wire \top/processor/sha_core/n3518_163 ;
wire \top/processor/sha_core/n3518_164 ;
wire \top/processor/sha_core/n3518_165 ;
wire \top/processor/sha_core/n3890_126 ;
wire \top/processor/sha_core/n3890_127 ;
wire \top/processor/sha_core/n3518_166 ;
wire \top/processor/sha_core/n3518_167 ;
wire \top/processor/sha_core/n3518_168 ;
wire \top/processor/sha_core/n3890_128 ;
wire \top/processor/sha_core/n3890_129 ;
wire \top/processor/sha_core/n3518_169 ;
wire \top/processor/sha_core/n3518_170 ;
wire \top/processor/sha_core/n3518_171 ;
wire \top/processor/sha_core/n3890_130 ;
wire \top/processor/sha_core/n3890_131 ;
wire \top/processor/sha_core/n3519_148 ;
wire \top/processor/sha_core/n3519_149 ;
wire \top/processor/sha_core/n3519_150 ;
wire \top/processor/sha_core/n3891_116 ;
wire \top/processor/sha_core/n3891_117 ;
wire \top/processor/sha_core/n3519_151 ;
wire \top/processor/sha_core/n3519_152 ;
wire \top/processor/sha_core/n3519_153 ;
wire \top/processor/sha_core/n3891_118 ;
wire \top/processor/sha_core/n3891_119 ;
wire \top/processor/sha_core/n3491_148 ;
wire \top/processor/sha_core/n3491_149 ;
wire \top/processor/sha_core/n3491_150 ;
wire \top/processor/sha_core/n3863_116 ;
wire \top/processor/sha_core/n3863_117 ;
wire \top/processor/sha_core/n3519_154 ;
wire \top/processor/sha_core/n3519_155 ;
wire \top/processor/sha_core/n3519_156 ;
wire \top/processor/sha_core/n3891_120 ;
wire \top/processor/sha_core/n3891_121 ;
wire \top/processor/sha_core/n3519_157 ;
wire \top/processor/sha_core/n3519_158 ;
wire \top/processor/sha_core/n3519_159 ;
wire \top/processor/sha_core/n3891_122 ;
wire \top/processor/sha_core/n3891_123 ;
wire \top/processor/sha_core/n3519_160 ;
wire \top/processor/sha_core/n3519_161 ;
wire \top/processor/sha_core/n3519_162 ;
wire \top/processor/sha_core/n3891_124 ;
wire \top/processor/sha_core/n3891_125 ;
wire \top/processor/sha_core/n3519_163 ;
wire \top/processor/sha_core/n3519_164 ;
wire \top/processor/sha_core/n3519_165 ;
wire \top/processor/sha_core/n3891_126 ;
wire \top/processor/sha_core/n3891_127 ;
wire \top/processor/sha_core/n3519_166 ;
wire \top/processor/sha_core/n3519_167 ;
wire \top/processor/sha_core/n3519_168 ;
wire \top/processor/sha_core/n3891_128 ;
wire \top/processor/sha_core/n3891_129 ;
wire \top/processor/sha_core/n3519_169 ;
wire \top/processor/sha_core/n3519_170 ;
wire \top/processor/sha_core/n3519_171 ;
wire \top/processor/sha_core/n3891_130 ;
wire \top/processor/sha_core/n3891_131 ;
wire \top/processor/sha_core/n3607_172 ;
wire \top/processor/sha_core/n3608_172 ;
wire \top/processor/sha_core/n3609_172 ;
wire \top/processor/sha_core/n3610_172 ;
wire \top/processor/sha_core/n3611_172 ;
wire \top/processor/sha_core/n3612_172 ;
wire \top/processor/sha_core/n3613_172 ;
wire \top/processor/sha_core/n3491_151 ;
wire \top/processor/sha_core/n3491_152 ;
wire \top/processor/sha_core/n3491_153 ;
wire \top/processor/sha_core/n3863_118 ;
wire \top/processor/sha_core/n3863_119 ;
wire \top/processor/sha_core/n3614_172 ;
wire \top/processor/sha_core/n3615_172 ;
wire \top/processor/sha_core/n3616_172 ;
wire \top/processor/sha_core/n3617_172 ;
wire \top/processor/sha_core/n3618_172 ;
wire \top/processor/sha_core/n3619_172 ;
wire \top/processor/sha_core/n3620_172 ;
wire \top/processor/sha_core/n3621_172 ;
wire \top/processor/sha_core/n3622_172 ;
wire \top/processor/sha_core/n3623_172 ;
wire \top/processor/sha_core/n3624_172 ;
wire \top/processor/sha_core/n3625_172 ;
wire \top/processor/sha_core/n3626_172 ;
wire \top/processor/sha_core/n3627_172 ;
wire \top/processor/sha_core/n3628_172 ;
wire \top/processor/sha_core/n3629_172 ;
wire \top/processor/sha_core/n3630_172 ;
wire \top/processor/sha_core/n3631_172 ;
wire \top/processor/sha_core/n3632_172 ;
wire \top/processor/sha_core/n3633_172 ;
wire \top/processor/sha_core/n3491_154 ;
wire \top/processor/sha_core/n3491_155 ;
wire \top/processor/sha_core/n3491_156 ;
wire \top/processor/sha_core/n3863_120 ;
wire \top/processor/sha_core/n3863_121 ;
wire \top/processor/sha_core/n3634_172 ;
wire \top/processor/sha_core/n3635_172 ;
wire \top/processor/sha_core/n3636_172 ;
wire \top/processor/sha_core/n3637_172 ;
wire \top/processor/sha_core/n3638_172 ;
wire \top/processor/sha_core/n3491_157 ;
wire \top/processor/sha_core/n3491_158 ;
wire \top/processor/sha_core/n3491_159 ;
wire \top/processor/sha_core/n3863_122 ;
wire \top/processor/sha_core/n3863_123 ;
wire \top/processor/sha_core/n3607_173 ;
wire \top/processor/sha_core/n3608_173 ;
wire \top/processor/sha_core/n3609_173 ;
wire \top/processor/sha_core/n3491_160 ;
wire \top/processor/sha_core/n3491_161 ;
wire \top/processor/sha_core/n3491_162 ;
wire \top/processor/sha_core/n3863_124 ;
wire \top/processor/sha_core/n3863_125 ;
wire \top/processor/sha_core/n3610_173 ;
wire \top/processor/sha_core/n3611_173 ;
wire \top/processor/sha_core/n3612_173 ;
wire \top/processor/sha_core/n3613_173 ;
wire \top/processor/sha_core/n3614_173 ;
wire \top/processor/sha_core/n3615_173 ;
wire \top/processor/sha_core/n3616_173 ;
wire \top/processor/sha_core/n3617_173 ;
wire \top/processor/sha_core/n3618_173 ;
wire \top/processor/sha_core/n3619_173 ;
wire \top/processor/sha_core/n3620_173 ;
wire \top/processor/sha_core/n3621_173 ;
wire \top/processor/sha_core/n3622_173 ;
wire \top/processor/sha_core/n3623_173 ;
wire \top/processor/sha_core/n3624_173 ;
wire \top/processor/sha_core/n3625_173 ;
wire \top/processor/sha_core/n3626_173 ;
wire \top/processor/sha_core/n3627_173 ;
wire \top/processor/sha_core/n3628_173 ;
wire \top/processor/sha_core/n3629_173 ;
wire \top/processor/sha_core/n3491_163 ;
wire \top/processor/sha_core/n3491_164 ;
wire \top/processor/sha_core/n3491_165 ;
wire \top/processor/sha_core/n3863_126 ;
wire \top/processor/sha_core/n3863_127 ;
wire \top/processor/sha_core/n3488_163 ;
wire \top/processor/sha_core/n3488_164 ;
wire \top/processor/sha_core/n3488_165 ;
wire \top/processor/sha_core/n3860_126 ;
wire \top/processor/sha_core/n3860_127 ;
wire \top/processor/sha_core/n3630_173 ;
wire \top/processor/sha_core/n3631_173 ;
wire \top/processor/sha_core/n3632_173 ;
wire \top/processor/sha_core/n3633_173 ;
wire \top/processor/sha_core/n3634_173 ;
wire \top/processor/sha_core/n3635_173 ;
wire \top/processor/sha_core/n3636_173 ;
wire \top/processor/sha_core/n3637_173 ;
wire \top/processor/sha_core/n3638_173 ;
wire \top/processor/sha_core/n3491_166 ;
wire \top/processor/sha_core/n3491_167 ;
wire \top/processor/sha_core/n3491_168 ;
wire \top/processor/sha_core/n3863_128 ;
wire \top/processor/sha_core/n3863_129 ;
wire \top/processor/sha_core/n3491_169 ;
wire \top/processor/sha_core/n3491_170 ;
wire \top/processor/sha_core/n3491_171 ;
wire \top/processor/sha_core/n3863_130 ;
wire \top/processor/sha_core/n3863_131 ;
wire \top/processor/sha_core/n3607_174 ;
wire \top/processor/sha_core/n3608_174 ;
wire \top/processor/sha_core/n3609_174 ;
wire \top/processor/sha_core/n3610_174 ;
wire \top/processor/sha_core/n3611_174 ;
wire \top/processor/sha_core/n3612_174 ;
wire \top/processor/sha_core/n3613_174 ;
wire \top/processor/sha_core/n3614_174 ;
wire \top/processor/sha_core/n3615_174 ;
wire \top/processor/sha_core/n3616_174 ;
wire \top/processor/sha_core/n3617_174 ;
wire \top/processor/sha_core/n3618_174 ;
wire \top/processor/sha_core/n3619_174 ;
wire \top/processor/sha_core/n3620_174 ;
wire \top/processor/sha_core/n3621_174 ;
wire \top/processor/sha_core/n3622_174 ;
wire \top/processor/sha_core/n3623_174 ;
wire \top/processor/sha_core/n3624_174 ;
wire \top/processor/sha_core/n3625_174 ;
wire \top/processor/sha_core/n3492_148 ;
wire \top/processor/sha_core/n3492_149 ;
wire \top/processor/sha_core/n3492_150 ;
wire \top/processor/sha_core/n3864_116 ;
wire \top/processor/sha_core/n3864_117 ;
wire \top/processor/sha_core/n3626_174 ;
wire \top/processor/sha_core/n3627_174 ;
wire \top/processor/sha_core/n3628_174 ;
wire \top/processor/sha_core/n3629_174 ;
wire \top/processor/sha_core/n3630_174 ;
wire \top/processor/sha_core/n3631_174 ;
wire \top/processor/sha_core/n3632_174 ;
wire \top/processor/sha_core/n3633_174 ;
wire \top/processor/sha_core/n3634_174 ;
wire \top/processor/sha_core/n3635_174 ;
wire \top/processor/sha_core/n3636_174 ;
wire \top/processor/sha_core/n3637_174 ;
wire \top/processor/sha_core/n3638_174 ;
wire \top/processor/sha_core/n3492_151 ;
wire \top/processor/sha_core/n3492_152 ;
wire \top/processor/sha_core/n3492_153 ;
wire \top/processor/sha_core/n3864_118 ;
wire \top/processor/sha_core/n3864_119 ;
wire \top/processor/sha_core/n3492_154 ;
wire \top/processor/sha_core/n3492_155 ;
wire \top/processor/sha_core/n3492_156 ;
wire \top/processor/sha_core/n3864_120 ;
wire \top/processor/sha_core/n3864_121 ;
wire \top/processor/sha_core/n3607_175 ;
wire \top/processor/sha_core/n3608_175 ;
wire \top/processor/sha_core/n3609_175 ;
wire \top/processor/sha_core/n3610_175 ;
wire \top/processor/sha_core/n3611_175 ;
wire \top/processor/sha_core/n3612_175 ;
wire \top/processor/sha_core/n3613_175 ;
wire \top/processor/sha_core/n3614_175 ;
wire \top/processor/sha_core/n3615_175 ;
wire \top/processor/sha_core/n3616_175 ;
wire \top/processor/sha_core/n3617_175 ;
wire \top/processor/sha_core/n3618_175 ;
wire \top/processor/sha_core/n3619_175 ;
wire \top/processor/sha_core/n3620_175 ;
wire \top/processor/sha_core/n3621_175 ;
wire \top/processor/sha_core/n3492_157 ;
wire \top/processor/sha_core/n3492_158 ;
wire \top/processor/sha_core/n3492_159 ;
wire \top/processor/sha_core/n3864_122 ;
wire \top/processor/sha_core/n3864_123 ;
wire \top/processor/sha_core/n3622_175 ;
wire \top/processor/sha_core/n3623_175 ;
wire \top/processor/sha_core/n3624_175 ;
wire \top/processor/sha_core/n3625_175 ;
wire \top/processor/sha_core/n3626_175 ;
wire \top/processor/sha_core/n3627_175 ;
wire \top/processor/sha_core/n3628_175 ;
wire \top/processor/sha_core/n3629_175 ;
wire \top/processor/sha_core/n3630_175 ;
wire \top/processor/sha_core/n3631_175 ;
wire \top/processor/sha_core/n3632_175 ;
wire \top/processor/sha_core/n3633_175 ;
wire \top/processor/sha_core/n3634_175 ;
wire \top/processor/sha_core/n3635_175 ;
wire \top/processor/sha_core/n3636_175 ;
wire \top/processor/sha_core/n3637_175 ;
wire \top/processor/sha_core/n3638_175 ;
wire \top/processor/sha_core/n3492_160 ;
wire \top/processor/sha_core/n3492_161 ;
wire \top/processor/sha_core/n3492_162 ;
wire \top/processor/sha_core/n3864_124 ;
wire \top/processor/sha_core/n3864_125 ;
wire \top/processor/sha_core/n3492_163 ;
wire \top/processor/sha_core/n3492_164 ;
wire \top/processor/sha_core/n3492_165 ;
wire \top/processor/sha_core/n3864_126 ;
wire \top/processor/sha_core/n3864_127 ;
wire \top/processor/sha_core/n3607_176 ;
wire \top/processor/sha_core/n3608_176 ;
wire \top/processor/sha_core/n3609_176 ;
wire \top/processor/sha_core/n3610_176 ;
wire \top/processor/sha_core/n3611_176 ;
wire \top/processor/sha_core/n3612_176 ;
wire \top/processor/sha_core/n3613_176 ;
wire \top/processor/sha_core/n3614_176 ;
wire \top/processor/sha_core/n3615_176 ;
wire \top/processor/sha_core/n3616_176 ;
wire \top/processor/sha_core/n3617_176 ;
wire \top/processor/sha_core/n3492_166 ;
wire \top/processor/sha_core/n3492_167 ;
wire \top/processor/sha_core/n3492_168 ;
wire \top/processor/sha_core/n3864_128 ;
wire \top/processor/sha_core/n3864_129 ;
wire \top/processor/sha_core/n3618_176 ;
wire \top/processor/sha_core/n3619_176 ;
wire \top/processor/sha_core/n3620_176 ;
wire \top/processor/sha_core/n3621_176 ;
wire \top/processor/sha_core/n3622_176 ;
wire \top/processor/sha_core/n3623_176 ;
wire \top/processor/sha_core/n3624_176 ;
wire \top/processor/sha_core/n3625_176 ;
wire \top/processor/sha_core/n3626_176 ;
wire \top/processor/sha_core/n3627_176 ;
wire \top/processor/sha_core/n3628_176 ;
wire \top/processor/sha_core/n3629_176 ;
wire \top/processor/sha_core/n3630_176 ;
wire \top/processor/sha_core/n3631_176 ;
wire \top/processor/sha_core/n3632_176 ;
wire \top/processor/sha_core/n3633_176 ;
wire \top/processor/sha_core/n3634_176 ;
wire \top/processor/sha_core/n3635_176 ;
wire \top/processor/sha_core/n3636_176 ;
wire \top/processor/sha_core/n3637_176 ;
wire \top/processor/sha_core/n3492_169 ;
wire \top/processor/sha_core/n3492_170 ;
wire \top/processor/sha_core/n3492_171 ;
wire \top/processor/sha_core/n3864_130 ;
wire \top/processor/sha_core/n3864_131 ;
wire \top/processor/sha_core/n3488_166 ;
wire \top/processor/sha_core/n3488_167 ;
wire \top/processor/sha_core/n3488_168 ;
wire \top/processor/sha_core/n3860_128 ;
wire \top/processor/sha_core/n3860_129 ;
wire \top/processor/sha_core/n3638_176 ;
wire \top/processor/sha_core/n3493_148 ;
wire \top/processor/sha_core/n3493_149 ;
wire \top/processor/sha_core/n3493_150 ;
wire \top/processor/sha_core/n3865_116 ;
wire \top/processor/sha_core/n3865_117 ;
wire \top/processor/sha_core/n3607_177 ;
wire \top/processor/sha_core/n3608_177 ;
wire \top/processor/sha_core/n3609_177 ;
wire \top/processor/sha_core/n3610_177 ;
wire \top/processor/sha_core/n3611_177 ;
wire \top/processor/sha_core/n3612_177 ;
wire \top/processor/sha_core/n3613_177 ;
wire \top/processor/sha_core/n3493_151 ;
wire \top/processor/sha_core/n3493_152 ;
wire \top/processor/sha_core/n3493_153 ;
wire \top/processor/sha_core/n3865_118 ;
wire \top/processor/sha_core/n3865_119 ;
wire \top/processor/sha_core/n3614_177 ;
wire \top/processor/sha_core/n3615_177 ;
wire \top/processor/sha_core/n3616_177 ;
wire \top/processor/sha_core/n3617_177 ;
wire \top/processor/sha_core/n3618_177 ;
wire \top/processor/sha_core/n3619_177 ;
wire \top/processor/sha_core/n3620_177 ;
wire \top/processor/sha_core/n3621_177 ;
wire \top/processor/sha_core/n3622_177 ;
wire \top/processor/sha_core/n3623_177 ;
wire \top/processor/sha_core/n3624_177 ;
wire \top/processor/sha_core/n3625_177 ;
wire \top/processor/sha_core/n3626_177 ;
wire \top/processor/sha_core/n3627_177 ;
wire \top/processor/sha_core/n3628_177 ;
wire \top/processor/sha_core/n3629_177 ;
wire \top/processor/sha_core/n3630_177 ;
wire \top/processor/sha_core/n3631_177 ;
wire \top/processor/sha_core/n3632_177 ;
wire \top/processor/sha_core/n3633_177 ;
wire \top/processor/sha_core/n3493_154 ;
wire \top/processor/sha_core/n3493_155 ;
wire \top/processor/sha_core/n3493_156 ;
wire \top/processor/sha_core/n3865_120 ;
wire \top/processor/sha_core/n3865_121 ;
wire \top/processor/sha_core/n3634_177 ;
wire \top/processor/sha_core/n3635_177 ;
wire \top/processor/sha_core/n3636_177 ;
wire \top/processor/sha_core/n3637_177 ;
wire \top/processor/sha_core/n3638_177 ;
wire \top/processor/sha_core/n3493_157 ;
wire \top/processor/sha_core/n3493_158 ;
wire \top/processor/sha_core/n3493_159 ;
wire \top/processor/sha_core/n3865_122 ;
wire \top/processor/sha_core/n3865_123 ;
wire \top/processor/sha_core/n3607_178 ;
wire \top/processor/sha_core/n3608_178 ;
wire \top/processor/sha_core/n3609_178 ;
wire \top/processor/sha_core/n3493_160 ;
wire \top/processor/sha_core/n3493_161 ;
wire \top/processor/sha_core/n3493_162 ;
wire \top/processor/sha_core/n3865_124 ;
wire \top/processor/sha_core/n3865_125 ;
wire \top/processor/sha_core/n3610_178 ;
wire \top/processor/sha_core/n3611_178 ;
wire \top/processor/sha_core/n3612_178 ;
wire \top/processor/sha_core/n3613_178 ;
wire \top/processor/sha_core/n3614_178 ;
wire \top/processor/sha_core/n3615_178 ;
wire \top/processor/sha_core/n3616_178 ;
wire \top/processor/sha_core/n3617_178 ;
wire \top/processor/sha_core/n3618_178 ;
wire \top/processor/sha_core/n3619_178 ;
wire \top/processor/sha_core/n3620_178 ;
wire \top/processor/sha_core/n3621_178 ;
wire \top/processor/sha_core/n3622_178 ;
wire \top/processor/sha_core/n3623_178 ;
wire \top/processor/sha_core/n3624_178 ;
wire \top/processor/sha_core/n3625_178 ;
wire \top/processor/sha_core/n3626_178 ;
wire \top/processor/sha_core/n3627_178 ;
wire \top/processor/sha_core/n3628_178 ;
wire \top/processor/sha_core/n3629_178 ;
wire \top/processor/sha_core/n3493_163 ;
wire \top/processor/sha_core/n3493_164 ;
wire \top/processor/sha_core/n3493_165 ;
wire \top/processor/sha_core/n3865_126 ;
wire \top/processor/sha_core/n3865_127 ;
wire \top/processor/sha_core/n3630_178 ;
wire \top/processor/sha_core/n3631_178 ;
wire \top/processor/sha_core/n3632_178 ;
wire \top/processor/sha_core/n3633_178 ;
wire \top/processor/sha_core/n3634_178 ;
wire \top/processor/sha_core/n3635_178 ;
wire \top/processor/sha_core/n3636_178 ;
wire \top/processor/sha_core/n3637_178 ;
wire \top/processor/sha_core/n3638_178 ;
wire \top/processor/sha_core/n3493_166 ;
wire \top/processor/sha_core/n3493_167 ;
wire \top/processor/sha_core/n3493_168 ;
wire \top/processor/sha_core/n3865_128 ;
wire \top/processor/sha_core/n3865_129 ;
wire \top/processor/sha_core/n3493_169 ;
wire \top/processor/sha_core/n3493_170 ;
wire \top/processor/sha_core/n3493_171 ;
wire \top/processor/sha_core/n3865_130 ;
wire \top/processor/sha_core/n3865_131 ;
wire \top/processor/sha_core/n3607_179 ;
wire \top/processor/sha_core/n3608_179 ;
wire \top/processor/sha_core/n3609_179 ;
wire \top/processor/sha_core/n3610_179 ;
wire \top/processor/sha_core/n3611_179 ;
wire \top/processor/sha_core/n3612_179 ;
wire \top/processor/sha_core/n3613_179 ;
wire \top/processor/sha_core/n3614_179 ;
wire \top/processor/sha_core/n3615_179 ;
wire \top/processor/sha_core/n3616_179 ;
wire \top/processor/sha_core/n3617_179 ;
wire \top/processor/sha_core/n3618_179 ;
wire \top/processor/sha_core/n3619_179 ;
wire \top/processor/sha_core/n3620_179 ;
wire \top/processor/sha_core/n3621_179 ;
wire \top/processor/sha_core/n3622_179 ;
wire \top/processor/sha_core/n3623_179 ;
wire \top/processor/sha_core/n3624_179 ;
wire \top/processor/sha_core/n3625_179 ;
wire \top/processor/sha_core/n3494_167 ;
wire \top/processor/sha_core/n3494_168 ;
wire \top/processor/sha_core/n3494_169 ;
wire \top/processor/sha_core/n3866_128 ;
wire \top/processor/sha_core/n3866_129 ;
wire \top/processor/sha_core/n3626_179 ;
wire \top/processor/sha_core/n3627_179 ;
wire \top/processor/sha_core/n3628_179 ;
wire \top/processor/sha_core/n3629_179 ;
wire \top/processor/sha_core/n3630_179 ;
wire \top/processor/sha_core/n3631_179 ;
wire \top/processor/sha_core/n3632_179 ;
wire \top/processor/sha_core/n3633_179 ;
wire \top/processor/sha_core/n3634_179 ;
wire \top/processor/sha_core/n3635_179 ;
wire \top/processor/sha_core/n3636_179 ;
wire \top/processor/sha_core/n3637_179 ;
wire \top/processor/sha_core/n3638_179 ;
wire \top/processor/sha_core/n3494_170 ;
wire \top/processor/sha_core/n3494_171 ;
wire \top/processor/sha_core/n3494_172 ;
wire \top/processor/sha_core/n3866_130 ;
wire \top/processor/sha_core/n3866_131 ;
wire \top/processor/sha_core/n3488_169 ;
wire \top/processor/sha_core/n3488_170 ;
wire \top/processor/sha_core/n3488_171 ;
wire \top/processor/sha_core/n3860_130 ;
wire \top/processor/sha_core/n3860_131 ;
wire \top/processor/sha_core/n3494_173 ;
wire \top/processor/sha_core/n3494_174 ;
wire \top/processor/sha_core/n3494_175 ;
wire \top/processor/sha_core/n3494_176 ;
wire \top/processor/sha_core/n3494_177 ;
wire \top/processor/sha_core/n3494_178 ;
wire \top/processor/sha_core/n3495_172 ;
wire \top/processor/sha_core/n3495_173 ;
wire \top/processor/sha_core/n3495_174 ;
wire \top/processor/sha_core/n3495_175 ;
wire \top/processor/sha_core/n3488_172 ;
wire \top/processor/sha_core/n3495_176 ;
wire \top/processor/sha_core/n3495_177 ;
wire \top/processor/sha_core/n3495_178 ;
wire \top/processor/sha_core/n3495_179 ;
wire \top/processor/sha_core/n3496_172 ;
wire \top/processor/sha_core/n3496_173 ;
wire \top/processor/sha_core/n3496_174 ;
wire \top/processor/sha_core/n3496_175 ;
wire \top/processor/sha_core/n3496_176 ;
wire \top/processor/sha_core/n3496_177 ;
wire \top/processor/sha_core/n3488_173 ;
wire \top/processor/sha_core/n3496_178 ;
wire \top/processor/sha_core/n3496_179 ;
wire \top/processor/sha_core/n3497_172 ;
wire \top/processor/sha_core/n3497_173 ;
wire \top/processor/sha_core/n3497_174 ;
wire \top/processor/sha_core/n3497_175 ;
wire \top/processor/sha_core/n3497_176 ;
wire \top/processor/sha_core/n3497_177 ;
wire \top/processor/sha_core/n3497_178 ;
wire \top/processor/sha_core/n3497_179 ;
wire \top/processor/sha_core/n3488_174 ;
wire \top/processor/sha_core/n3498_172 ;
wire \top/processor/sha_core/n3498_173 ;
wire \top/processor/sha_core/n3498_174 ;
wire \top/processor/sha_core/n3498_175 ;
wire \top/processor/sha_core/n3498_176 ;
wire \top/processor/sha_core/n3498_177 ;
wire \top/processor/sha_core/n3498_178 ;
wire \top/processor/sha_core/n3498_179 ;
wire \top/processor/sha_core/n3499_172 ;
wire \top/processor/sha_core/n3499_173 ;
wire \top/processor/sha_core/n3489_172 ;
wire \top/processor/sha_core/n3499_174 ;
wire \top/processor/sha_core/n3499_175 ;
wire \top/processor/sha_core/n3499_176 ;
wire \top/processor/sha_core/n3499_177 ;
wire \top/processor/sha_core/n3499_178 ;
wire \top/processor/sha_core/n3499_179 ;
wire \top/processor/sha_core/n3500_172 ;
wire \top/processor/sha_core/n3500_173 ;
wire \top/processor/sha_core/n3500_174 ;
wire \top/processor/sha_core/n3500_175 ;
wire \top/processor/sha_core/n3489_173 ;
wire \top/processor/sha_core/n3488_175 ;
wire \top/processor/sha_core/n3500_176 ;
wire \top/processor/sha_core/n3500_177 ;
wire \top/processor/sha_core/n3500_178 ;
wire \top/processor/sha_core/n3500_179 ;
wire \top/processor/sha_core/n3501_172 ;
wire \top/processor/sha_core/n3501_173 ;
wire \top/processor/sha_core/n3501_174 ;
wire \top/processor/sha_core/n3501_175 ;
wire \top/processor/sha_core/n3501_176 ;
wire \top/processor/sha_core/n3501_177 ;
wire \top/processor/sha_core/n3489_174 ;
wire \top/processor/sha_core/n3501_178 ;
wire \top/processor/sha_core/n3501_179 ;
wire \top/processor/sha_core/n3502_172 ;
wire \top/processor/sha_core/n3502_173 ;
wire \top/processor/sha_core/n3502_174 ;
wire \top/processor/sha_core/n3502_175 ;
wire \top/processor/sha_core/n3502_176 ;
wire \top/processor/sha_core/n3502_177 ;
wire \top/processor/sha_core/n3502_178 ;
wire \top/processor/sha_core/n3502_179 ;
wire \top/processor/sha_core/n3489_175 ;
wire \top/processor/sha_core/n3503_172 ;
wire \top/processor/sha_core/n3503_173 ;
wire \top/processor/sha_core/n3503_174 ;
wire \top/processor/sha_core/n3503_175 ;
wire \top/processor/sha_core/n3503_176 ;
wire \top/processor/sha_core/n3503_177 ;
wire \top/processor/sha_core/n3503_178 ;
wire \top/processor/sha_core/n3503_179 ;
wire \top/processor/sha_core/n3504_172 ;
wire \top/processor/sha_core/n3504_173 ;
wire \top/processor/sha_core/n3489_176 ;
wire \top/processor/sha_core/n3504_174 ;
wire \top/processor/sha_core/n3504_175 ;
wire \top/processor/sha_core/n3504_176 ;
wire \top/processor/sha_core/n3504_177 ;
wire \top/processor/sha_core/n3504_178 ;
wire \top/processor/sha_core/n3504_179 ;
wire \top/processor/sha_core/n3505_172 ;
wire \top/processor/sha_core/n3505_173 ;
wire \top/processor/sha_core/n3505_174 ;
wire \top/processor/sha_core/n3505_175 ;
wire \top/processor/sha_core/n3489_177 ;
wire \top/processor/sha_core/n3505_176 ;
wire \top/processor/sha_core/n3505_177 ;
wire \top/processor/sha_core/n3505_178 ;
wire \top/processor/sha_core/n3505_179 ;
wire \top/processor/sha_core/n3506_172 ;
wire \top/processor/sha_core/n3506_173 ;
wire \top/processor/sha_core/n3506_174 ;
wire \top/processor/sha_core/n3506_175 ;
wire \top/processor/sha_core/n3506_176 ;
wire \top/processor/sha_core/n3506_177 ;
wire \top/processor/sha_core/n3489_178 ;
wire \top/processor/sha_core/n3506_178 ;
wire \top/processor/sha_core/n3506_179 ;
wire \top/processor/sha_core/n3507_172 ;
wire \top/processor/sha_core/n3507_173 ;
wire \top/processor/sha_core/n3507_174 ;
wire \top/processor/sha_core/n3507_175 ;
wire \top/processor/sha_core/n3507_176 ;
wire \top/processor/sha_core/n3507_177 ;
wire \top/processor/sha_core/n3507_178 ;
wire \top/processor/sha_core/n3507_179 ;
wire \top/processor/sha_core/n3489_179 ;
wire \top/processor/sha_core/n3508_172 ;
wire \top/processor/sha_core/n3508_173 ;
wire \top/processor/sha_core/n3508_174 ;
wire \top/processor/sha_core/n3508_175 ;
wire \top/processor/sha_core/n3508_176 ;
wire \top/processor/sha_core/n3508_177 ;
wire \top/processor/sha_core/n3508_178 ;
wire \top/processor/sha_core/n3508_179 ;
wire \top/processor/sha_core/n3509_172 ;
wire \top/processor/sha_core/n3509_173 ;
wire \top/processor/sha_core/n3490_172 ;
wire \top/processor/sha_core/n3509_174 ;
wire \top/processor/sha_core/n3509_175 ;
wire \top/processor/sha_core/n3509_176 ;
wire \top/processor/sha_core/n3509_177 ;
wire \top/processor/sha_core/n3509_178 ;
wire \top/processor/sha_core/n3509_179 ;
wire \top/processor/sha_core/n3510_172 ;
wire \top/processor/sha_core/n3510_173 ;
wire \top/processor/sha_core/n3510_174 ;
wire \top/processor/sha_core/n3510_175 ;
wire \top/processor/sha_core/n3490_173 ;
wire \top/processor/sha_core/n3510_176 ;
wire \top/processor/sha_core/n3510_177 ;
wire \top/processor/sha_core/n3510_178 ;
wire \top/processor/sha_core/n3510_179 ;
wire \top/processor/sha_core/n3511_172 ;
wire \top/processor/sha_core/n3511_173 ;
wire \top/processor/sha_core/n3511_174 ;
wire \top/processor/sha_core/n3511_175 ;
wire \top/processor/sha_core/n3511_176 ;
wire \top/processor/sha_core/n3511_177 ;
wire \top/processor/sha_core/n3490_174 ;
wire \top/processor/sha_core/n3511_178 ;
wire \top/processor/sha_core/n3511_179 ;
wire \top/processor/sha_core/n3512_172 ;
wire \top/processor/sha_core/n3512_173 ;
wire \top/processor/sha_core/n3512_174 ;
wire \top/processor/sha_core/n3512_175 ;
wire \top/processor/sha_core/n3512_176 ;
wire \top/processor/sha_core/n3512_177 ;
wire \top/processor/sha_core/n3512_178 ;
wire \top/processor/sha_core/n3512_179 ;
wire \top/processor/sha_core/n3490_175 ;
wire \top/processor/sha_core/n3488_176 ;
wire \top/processor/sha_core/n3513_172 ;
wire \top/processor/sha_core/n3513_173 ;
wire \top/processor/sha_core/n3513_174 ;
wire \top/processor/sha_core/n3513_175 ;
wire \top/processor/sha_core/n3513_176 ;
wire \top/processor/sha_core/n3513_177 ;
wire \top/processor/sha_core/n3513_178 ;
wire \top/processor/sha_core/n3513_179 ;
wire \top/processor/sha_core/n3514_172 ;
wire \top/processor/sha_core/n3514_173 ;
wire \top/processor/sha_core/n3490_176 ;
wire \top/processor/sha_core/n3514_174 ;
wire \top/processor/sha_core/n3514_175 ;
wire \top/processor/sha_core/n3514_176 ;
wire \top/processor/sha_core/n3514_177 ;
wire \top/processor/sha_core/n3514_178 ;
wire \top/processor/sha_core/n3514_179 ;
wire \top/processor/sha_core/n3515_172 ;
wire \top/processor/sha_core/n3515_173 ;
wire \top/processor/sha_core/n3515_174 ;
wire \top/processor/sha_core/n3515_175 ;
wire \top/processor/sha_core/n3490_177 ;
wire \top/processor/sha_core/n3515_176 ;
wire \top/processor/sha_core/n3515_177 ;
wire \top/processor/sha_core/n3515_178 ;
wire \top/processor/sha_core/n3515_179 ;
wire \top/processor/sha_core/n3516_172 ;
wire \top/processor/sha_core/n3516_173 ;
wire \top/processor/sha_core/n3516_174 ;
wire \top/processor/sha_core/n3516_175 ;
wire \top/processor/sha_core/n3516_176 ;
wire \top/processor/sha_core/n3516_177 ;
wire \top/processor/sha_core/n3490_178 ;
wire \top/processor/sha_core/n3516_178 ;
wire \top/processor/sha_core/n3516_179 ;
wire \top/processor/sha_core/n3517_172 ;
wire \top/processor/sha_core/n3517_173 ;
wire \top/processor/sha_core/n3517_174 ;
wire \top/processor/sha_core/n3517_175 ;
wire \top/processor/sha_core/n3517_176 ;
wire \top/processor/sha_core/n3517_177 ;
wire \top/processor/sha_core/n3517_178 ;
wire \top/processor/sha_core/n3517_179 ;
wire \top/processor/sha_core/n3490_179 ;
wire \top/processor/sha_core/n3518_172 ;
wire \top/processor/sha_core/n3518_173 ;
wire \top/processor/sha_core/n3518_174 ;
wire \top/processor/sha_core/n3518_175 ;
wire \top/processor/sha_core/n3518_176 ;
wire \top/processor/sha_core/n3518_177 ;
wire \top/processor/sha_core/n3518_178 ;
wire \top/processor/sha_core/n3518_179 ;
wire \top/processor/sha_core/n3519_172 ;
wire \top/processor/sha_core/n3519_173 ;
wire \top/processor/sha_core/n3491_172 ;
wire \top/processor/sha_core/n3519_174 ;
wire \top/processor/sha_core/n3519_175 ;
wire \top/processor/sha_core/n3519_176 ;
wire \top/processor/sha_core/n3519_177 ;
wire \top/processor/sha_core/n3519_178 ;
wire \top/processor/sha_core/n3519_179 ;
wire \top/processor/sha_core/n3491_173 ;
wire \top/processor/sha_core/n3491_174 ;
wire \top/processor/sha_core/n3491_175 ;
wire \top/processor/sha_core/n3491_176 ;
wire \top/processor/sha_core/n3491_177 ;
wire \top/processor/sha_core/n3488_177 ;
wire \top/processor/sha_core/n3491_178 ;
wire \top/processor/sha_core/n3491_179 ;
wire \top/processor/sha_core/n3492_172 ;
wire \top/processor/sha_core/n3492_173 ;
wire \top/processor/sha_core/n3492_174 ;
wire \top/processor/sha_core/n3492_175 ;
wire \top/processor/sha_core/n3492_176 ;
wire \top/processor/sha_core/n3492_177 ;
wire \top/processor/sha_core/n3492_178 ;
wire \top/processor/sha_core/n3492_179 ;
wire \top/processor/sha_core/n3488_178 ;
wire \top/processor/sha_core/n3493_172 ;
wire \top/processor/sha_core/n3493_173 ;
wire \top/processor/sha_core/n3493_174 ;
wire \top/processor/sha_core/n3493_175 ;
wire \top/processor/sha_core/n3493_176 ;
wire \top/processor/sha_core/n3493_177 ;
wire \top/processor/sha_core/n3493_178 ;
wire \top/processor/sha_core/n3493_179 ;
wire \top/processor/sha_core/n3494_179 ;
wire \top/processor/sha_core/n3494_180 ;
wire \top/processor/sha_core/n3488_179 ;
wire \top/processor/sha_core/n327_132 ;
wire \top/processor/sha_core/n327_133 ;
wire \top/processor/sha_core/n327_134 ;
wire \top/processor/sha_core/n327_135 ;
wire \top/processor/sha_core/n327_136 ;
wire \top/processor/sha_core/n327_137 ;
wire \top/processor/sha_core/n327_138 ;
wire \top/processor/sha_core/n327_139 ;
wire \top/processor/sha_core/n327_140 ;
wire \top/processor/sha_core/n327_141 ;
wire \top/processor/sha_core/n327_142 ;
wire \top/processor/sha_core/n327_143 ;
wire \top/processor/sha_core/n327_144 ;
wire \top/processor/sha_core/n327_145 ;
wire \top/processor/sha_core/n327_146 ;
wire \top/processor/sha_core/n327_147 ;
wire \top/processor/sha_core/n327_148 ;
wire \top/processor/sha_core/n327_149 ;
wire \top/processor/sha_core/n327_150 ;
wire \top/processor/sha_core/n327_151 ;
wire \top/processor/sha_core/n327_152 ;
wire \top/processor/sha_core/n327_153 ;
wire \top/processor/sha_core/n327_154 ;
wire \top/processor/sha_core/n327_155 ;
wire \top/processor/sha_core/n327_156 ;
wire \top/processor/sha_core/n327_157 ;
wire \top/processor/sha_core/n327_158 ;
wire \top/processor/sha_core/n327_159 ;
wire \top/processor/sha_core/n327_160 ;
wire \top/processor/sha_core/n327_161 ;
wire \top/processor/sha_core/n327_162 ;
wire \top/processor/sha_core/n327_163 ;
wire \top/processor/sha_core/n328_132 ;
wire \top/processor/sha_core/n328_133 ;
wire \top/processor/sha_core/n328_134 ;
wire \top/processor/sha_core/n328_135 ;
wire \top/processor/sha_core/n328_136 ;
wire \top/processor/sha_core/n328_137 ;
wire \top/processor/sha_core/n328_138 ;
wire \top/processor/sha_core/n328_139 ;
wire \top/processor/sha_core/n328_140 ;
wire \top/processor/sha_core/n328_141 ;
wire \top/processor/sha_core/n328_142 ;
wire \top/processor/sha_core/n328_143 ;
wire \top/processor/sha_core/n328_144 ;
wire \top/processor/sha_core/n328_145 ;
wire \top/processor/sha_core/n328_146 ;
wire \top/processor/sha_core/n328_147 ;
wire \top/processor/sha_core/n328_148 ;
wire \top/processor/sha_core/n328_149 ;
wire \top/processor/sha_core/n328_150 ;
wire \top/processor/sha_core/n328_151 ;
wire \top/processor/sha_core/n328_152 ;
wire \top/processor/sha_core/n328_153 ;
wire \top/processor/sha_core/n328_154 ;
wire \top/processor/sha_core/n328_155 ;
wire \top/processor/sha_core/n328_156 ;
wire \top/processor/sha_core/n328_157 ;
wire \top/processor/sha_core/n328_158 ;
wire \top/processor/sha_core/n328_159 ;
wire \top/processor/sha_core/n328_160 ;
wire \top/processor/sha_core/n328_161 ;
wire \top/processor/sha_core/n328_162 ;
wire \top/processor/sha_core/n328_163 ;
wire \top/processor/sha_core/n329_132 ;
wire \top/processor/sha_core/n329_133 ;
wire \top/processor/sha_core/n329_134 ;
wire \top/processor/sha_core/n329_135 ;
wire \top/processor/sha_core/n329_136 ;
wire \top/processor/sha_core/n329_137 ;
wire \top/processor/sha_core/n329_138 ;
wire \top/processor/sha_core/n329_139 ;
wire \top/processor/sha_core/n329_140 ;
wire \top/processor/sha_core/n329_141 ;
wire \top/processor/sha_core/n329_142 ;
wire \top/processor/sha_core/n329_143 ;
wire \top/processor/sha_core/n329_144 ;
wire \top/processor/sha_core/n329_145 ;
wire \top/processor/sha_core/n329_146 ;
wire \top/processor/sha_core/n329_147 ;
wire \top/processor/sha_core/n329_148 ;
wire \top/processor/sha_core/n329_149 ;
wire \top/processor/sha_core/n329_150 ;
wire \top/processor/sha_core/n329_151 ;
wire \top/processor/sha_core/n329_152 ;
wire \top/processor/sha_core/n329_153 ;
wire \top/processor/sha_core/n329_154 ;
wire \top/processor/sha_core/n329_155 ;
wire \top/processor/sha_core/n329_156 ;
wire \top/processor/sha_core/n329_157 ;
wire \top/processor/sha_core/n329_158 ;
wire \top/processor/sha_core/n329_159 ;
wire \top/processor/sha_core/n329_160 ;
wire \top/processor/sha_core/n329_161 ;
wire \top/processor/sha_core/n329_162 ;
wire \top/processor/sha_core/n329_163 ;
wire \top/processor/sha_core/n330_132 ;
wire \top/processor/sha_core/n330_133 ;
wire \top/processor/sha_core/n330_134 ;
wire \top/processor/sha_core/n330_135 ;
wire \top/processor/sha_core/n330_136 ;
wire \top/processor/sha_core/n330_137 ;
wire \top/processor/sha_core/n330_138 ;
wire \top/processor/sha_core/n330_139 ;
wire \top/processor/sha_core/n330_140 ;
wire \top/processor/sha_core/n330_141 ;
wire \top/processor/sha_core/n330_142 ;
wire \top/processor/sha_core/n330_143 ;
wire \top/processor/sha_core/n330_144 ;
wire \top/processor/sha_core/n330_145 ;
wire \top/processor/sha_core/n330_146 ;
wire \top/processor/sha_core/n330_147 ;
wire \top/processor/sha_core/n330_148 ;
wire \top/processor/sha_core/n330_149 ;
wire \top/processor/sha_core/n330_150 ;
wire \top/processor/sha_core/n330_151 ;
wire \top/processor/sha_core/n330_152 ;
wire \top/processor/sha_core/n330_153 ;
wire \top/processor/sha_core/n330_154 ;
wire \top/processor/sha_core/n330_155 ;
wire \top/processor/sha_core/n330_156 ;
wire \top/processor/sha_core/n330_157 ;
wire \top/processor/sha_core/n330_158 ;
wire \top/processor/sha_core/n330_159 ;
wire \top/processor/sha_core/n330_160 ;
wire \top/processor/sha_core/n330_161 ;
wire \top/processor/sha_core/n330_162 ;
wire \top/processor/sha_core/n330_163 ;
wire \top/processor/sha_core/n331_132 ;
wire \top/processor/sha_core/n331_133 ;
wire \top/processor/sha_core/n331_134 ;
wire \top/processor/sha_core/n331_135 ;
wire \top/processor/sha_core/n331_136 ;
wire \top/processor/sha_core/n331_137 ;
wire \top/processor/sha_core/n331_138 ;
wire \top/processor/sha_core/n331_139 ;
wire \top/processor/sha_core/n331_140 ;
wire \top/processor/sha_core/n331_141 ;
wire \top/processor/sha_core/n331_142 ;
wire \top/processor/sha_core/n331_143 ;
wire \top/processor/sha_core/n331_144 ;
wire \top/processor/sha_core/n331_145 ;
wire \top/processor/sha_core/n331_146 ;
wire \top/processor/sha_core/n331_147 ;
wire \top/processor/sha_core/n331_148 ;
wire \top/processor/sha_core/n331_149 ;
wire \top/processor/sha_core/n331_150 ;
wire \top/processor/sha_core/n331_151 ;
wire \top/processor/sha_core/n331_152 ;
wire \top/processor/sha_core/n331_153 ;
wire \top/processor/sha_core/n331_154 ;
wire \top/processor/sha_core/n331_155 ;
wire \top/processor/sha_core/n331_156 ;
wire \top/processor/sha_core/n331_157 ;
wire \top/processor/sha_core/n331_158 ;
wire \top/processor/sha_core/n331_159 ;
wire \top/processor/sha_core/n331_160 ;
wire \top/processor/sha_core/n331_161 ;
wire \top/processor/sha_core/n331_162 ;
wire \top/processor/sha_core/n331_163 ;
wire \top/processor/sha_core/n332_132 ;
wire \top/processor/sha_core/n332_133 ;
wire \top/processor/sha_core/n332_134 ;
wire \top/processor/sha_core/n332_135 ;
wire \top/processor/sha_core/n332_136 ;
wire \top/processor/sha_core/n332_137 ;
wire \top/processor/sha_core/n332_138 ;
wire \top/processor/sha_core/n332_139 ;
wire \top/processor/sha_core/n332_140 ;
wire \top/processor/sha_core/n332_141 ;
wire \top/processor/sha_core/n332_142 ;
wire \top/processor/sha_core/n332_143 ;
wire \top/processor/sha_core/n332_144 ;
wire \top/processor/sha_core/n332_145 ;
wire \top/processor/sha_core/n332_146 ;
wire \top/processor/sha_core/n332_147 ;
wire \top/processor/sha_core/n332_148 ;
wire \top/processor/sha_core/n332_149 ;
wire \top/processor/sha_core/n332_150 ;
wire \top/processor/sha_core/n332_151 ;
wire \top/processor/sha_core/n332_152 ;
wire \top/processor/sha_core/n332_153 ;
wire \top/processor/sha_core/n332_154 ;
wire \top/processor/sha_core/n332_155 ;
wire \top/processor/sha_core/n332_156 ;
wire \top/processor/sha_core/n332_157 ;
wire \top/processor/sha_core/n332_158 ;
wire \top/processor/sha_core/n332_159 ;
wire \top/processor/sha_core/n332_160 ;
wire \top/processor/sha_core/n332_161 ;
wire \top/processor/sha_core/n332_162 ;
wire \top/processor/sha_core/n332_163 ;
wire \top/processor/sha_core/n333_132 ;
wire \top/processor/sha_core/n333_133 ;
wire \top/processor/sha_core/n333_134 ;
wire \top/processor/sha_core/n333_135 ;
wire \top/processor/sha_core/n333_136 ;
wire \top/processor/sha_core/n333_137 ;
wire \top/processor/sha_core/n333_138 ;
wire \top/processor/sha_core/n333_139 ;
wire \top/processor/sha_core/n333_140 ;
wire \top/processor/sha_core/n333_141 ;
wire \top/processor/sha_core/n333_142 ;
wire \top/processor/sha_core/n333_143 ;
wire \top/processor/sha_core/n333_144 ;
wire \top/processor/sha_core/n333_145 ;
wire \top/processor/sha_core/n333_146 ;
wire \top/processor/sha_core/n333_147 ;
wire \top/processor/sha_core/n333_148 ;
wire \top/processor/sha_core/n333_149 ;
wire \top/processor/sha_core/n333_150 ;
wire \top/processor/sha_core/n333_151 ;
wire \top/processor/sha_core/n333_152 ;
wire \top/processor/sha_core/n333_153 ;
wire \top/processor/sha_core/n333_154 ;
wire \top/processor/sha_core/n333_155 ;
wire \top/processor/sha_core/n333_156 ;
wire \top/processor/sha_core/n333_157 ;
wire \top/processor/sha_core/n333_158 ;
wire \top/processor/sha_core/n333_159 ;
wire \top/processor/sha_core/n333_160 ;
wire \top/processor/sha_core/n333_161 ;
wire \top/processor/sha_core/n333_162 ;
wire \top/processor/sha_core/n333_163 ;
wire \top/processor/sha_core/n334_132 ;
wire \top/processor/sha_core/n334_133 ;
wire \top/processor/sha_core/n334_134 ;
wire \top/processor/sha_core/n334_135 ;
wire \top/processor/sha_core/n334_136 ;
wire \top/processor/sha_core/n334_137 ;
wire \top/processor/sha_core/n334_138 ;
wire \top/processor/sha_core/n334_139 ;
wire \top/processor/sha_core/n334_140 ;
wire \top/processor/sha_core/n334_141 ;
wire \top/processor/sha_core/n334_142 ;
wire \top/processor/sha_core/n334_143 ;
wire \top/processor/sha_core/n334_144 ;
wire \top/processor/sha_core/n334_145 ;
wire \top/processor/sha_core/n334_146 ;
wire \top/processor/sha_core/n334_147 ;
wire \top/processor/sha_core/n334_148 ;
wire \top/processor/sha_core/n334_149 ;
wire \top/processor/sha_core/n334_150 ;
wire \top/processor/sha_core/n334_151 ;
wire \top/processor/sha_core/n334_152 ;
wire \top/processor/sha_core/n334_153 ;
wire \top/processor/sha_core/n334_154 ;
wire \top/processor/sha_core/n334_155 ;
wire \top/processor/sha_core/n334_156 ;
wire \top/processor/sha_core/n334_157 ;
wire \top/processor/sha_core/n334_158 ;
wire \top/processor/sha_core/n334_159 ;
wire \top/processor/sha_core/n334_160 ;
wire \top/processor/sha_core/n334_161 ;
wire \top/processor/sha_core/n334_162 ;
wire \top/processor/sha_core/n334_163 ;
wire \top/processor/sha_core/n335_132 ;
wire \top/processor/sha_core/n335_133 ;
wire \top/processor/sha_core/n335_134 ;
wire \top/processor/sha_core/n335_135 ;
wire \top/processor/sha_core/n335_136 ;
wire \top/processor/sha_core/n335_137 ;
wire \top/processor/sha_core/n335_138 ;
wire \top/processor/sha_core/n335_139 ;
wire \top/processor/sha_core/n335_140 ;
wire \top/processor/sha_core/n335_141 ;
wire \top/processor/sha_core/n335_142 ;
wire \top/processor/sha_core/n335_143 ;
wire \top/processor/sha_core/n335_144 ;
wire \top/processor/sha_core/n335_145 ;
wire \top/processor/sha_core/n335_146 ;
wire \top/processor/sha_core/n335_147 ;
wire \top/processor/sha_core/n335_148 ;
wire \top/processor/sha_core/n335_149 ;
wire \top/processor/sha_core/n335_150 ;
wire \top/processor/sha_core/n335_151 ;
wire \top/processor/sha_core/n335_152 ;
wire \top/processor/sha_core/n335_153 ;
wire \top/processor/sha_core/n335_154 ;
wire \top/processor/sha_core/n335_155 ;
wire \top/processor/sha_core/n335_156 ;
wire \top/processor/sha_core/n335_157 ;
wire \top/processor/sha_core/n335_158 ;
wire \top/processor/sha_core/n335_159 ;
wire \top/processor/sha_core/n335_160 ;
wire \top/processor/sha_core/n335_161 ;
wire \top/processor/sha_core/n335_162 ;
wire \top/processor/sha_core/n335_163 ;
wire \top/processor/sha_core/n336_132 ;
wire \top/processor/sha_core/n336_133 ;
wire \top/processor/sha_core/n336_134 ;
wire \top/processor/sha_core/n336_135 ;
wire \top/processor/sha_core/n336_136 ;
wire \top/processor/sha_core/n336_137 ;
wire \top/processor/sha_core/n336_138 ;
wire \top/processor/sha_core/n336_139 ;
wire \top/processor/sha_core/n336_140 ;
wire \top/processor/sha_core/n336_141 ;
wire \top/processor/sha_core/n336_142 ;
wire \top/processor/sha_core/n336_143 ;
wire \top/processor/sha_core/n336_144 ;
wire \top/processor/sha_core/n336_145 ;
wire \top/processor/sha_core/n336_146 ;
wire \top/processor/sha_core/n336_147 ;
wire \top/processor/sha_core/n336_148 ;
wire \top/processor/sha_core/n336_149 ;
wire \top/processor/sha_core/n336_150 ;
wire \top/processor/sha_core/n336_151 ;
wire \top/processor/sha_core/n336_152 ;
wire \top/processor/sha_core/n336_153 ;
wire \top/processor/sha_core/n336_154 ;
wire \top/processor/sha_core/n336_155 ;
wire \top/processor/sha_core/n336_156 ;
wire \top/processor/sha_core/n336_157 ;
wire \top/processor/sha_core/n336_158 ;
wire \top/processor/sha_core/n336_159 ;
wire \top/processor/sha_core/n336_160 ;
wire \top/processor/sha_core/n336_161 ;
wire \top/processor/sha_core/n336_162 ;
wire \top/processor/sha_core/n336_163 ;
wire \top/processor/sha_core/n337_132 ;
wire \top/processor/sha_core/n337_133 ;
wire \top/processor/sha_core/n337_134 ;
wire \top/processor/sha_core/n337_135 ;
wire \top/processor/sha_core/n337_136 ;
wire \top/processor/sha_core/n337_137 ;
wire \top/processor/sha_core/n337_138 ;
wire \top/processor/sha_core/n337_139 ;
wire \top/processor/sha_core/n337_140 ;
wire \top/processor/sha_core/n337_141 ;
wire \top/processor/sha_core/n337_142 ;
wire \top/processor/sha_core/n337_143 ;
wire \top/processor/sha_core/n337_144 ;
wire \top/processor/sha_core/n337_145 ;
wire \top/processor/sha_core/n337_146 ;
wire \top/processor/sha_core/n337_147 ;
wire \top/processor/sha_core/n337_148 ;
wire \top/processor/sha_core/n337_149 ;
wire \top/processor/sha_core/n337_150 ;
wire \top/processor/sha_core/n337_151 ;
wire \top/processor/sha_core/n337_152 ;
wire \top/processor/sha_core/n337_153 ;
wire \top/processor/sha_core/n337_154 ;
wire \top/processor/sha_core/n337_155 ;
wire \top/processor/sha_core/n337_156 ;
wire \top/processor/sha_core/n337_157 ;
wire \top/processor/sha_core/n337_158 ;
wire \top/processor/sha_core/n337_159 ;
wire \top/processor/sha_core/n337_160 ;
wire \top/processor/sha_core/n337_161 ;
wire \top/processor/sha_core/n337_162 ;
wire \top/processor/sha_core/n337_163 ;
wire \top/processor/sha_core/n338_132 ;
wire \top/processor/sha_core/n338_133 ;
wire \top/processor/sha_core/n338_134 ;
wire \top/processor/sha_core/n338_135 ;
wire \top/processor/sha_core/n338_136 ;
wire \top/processor/sha_core/n338_137 ;
wire \top/processor/sha_core/n338_138 ;
wire \top/processor/sha_core/n338_139 ;
wire \top/processor/sha_core/n338_140 ;
wire \top/processor/sha_core/n338_141 ;
wire \top/processor/sha_core/n338_142 ;
wire \top/processor/sha_core/n338_143 ;
wire \top/processor/sha_core/n338_144 ;
wire \top/processor/sha_core/n338_145 ;
wire \top/processor/sha_core/n338_146 ;
wire \top/processor/sha_core/n338_147 ;
wire \top/processor/sha_core/n338_148 ;
wire \top/processor/sha_core/n338_149 ;
wire \top/processor/sha_core/n338_150 ;
wire \top/processor/sha_core/n338_151 ;
wire \top/processor/sha_core/n338_152 ;
wire \top/processor/sha_core/n338_153 ;
wire \top/processor/sha_core/n338_154 ;
wire \top/processor/sha_core/n338_155 ;
wire \top/processor/sha_core/n338_156 ;
wire \top/processor/sha_core/n338_157 ;
wire \top/processor/sha_core/n338_158 ;
wire \top/processor/sha_core/n338_159 ;
wire \top/processor/sha_core/n338_160 ;
wire \top/processor/sha_core/n338_161 ;
wire \top/processor/sha_core/n338_162 ;
wire \top/processor/sha_core/n338_163 ;
wire \top/processor/sha_core/n339_132 ;
wire \top/processor/sha_core/n339_133 ;
wire \top/processor/sha_core/n339_134 ;
wire \top/processor/sha_core/n339_135 ;
wire \top/processor/sha_core/n339_136 ;
wire \top/processor/sha_core/n339_137 ;
wire \top/processor/sha_core/n339_138 ;
wire \top/processor/sha_core/n339_139 ;
wire \top/processor/sha_core/n339_140 ;
wire \top/processor/sha_core/n339_141 ;
wire \top/processor/sha_core/n339_142 ;
wire \top/processor/sha_core/n339_143 ;
wire \top/processor/sha_core/n339_144 ;
wire \top/processor/sha_core/n339_145 ;
wire \top/processor/sha_core/n339_146 ;
wire \top/processor/sha_core/n339_147 ;
wire \top/processor/sha_core/n339_148 ;
wire \top/processor/sha_core/n339_149 ;
wire \top/processor/sha_core/n339_150 ;
wire \top/processor/sha_core/n339_151 ;
wire \top/processor/sha_core/n339_152 ;
wire \top/processor/sha_core/n339_153 ;
wire \top/processor/sha_core/n339_154 ;
wire \top/processor/sha_core/n339_155 ;
wire \top/processor/sha_core/n339_156 ;
wire \top/processor/sha_core/n339_157 ;
wire \top/processor/sha_core/n339_158 ;
wire \top/processor/sha_core/n339_159 ;
wire \top/processor/sha_core/n339_160 ;
wire \top/processor/sha_core/n339_161 ;
wire \top/processor/sha_core/n339_162 ;
wire \top/processor/sha_core/n339_163 ;
wire \top/processor/sha_core/n340_132 ;
wire \top/processor/sha_core/n340_133 ;
wire \top/processor/sha_core/n340_134 ;
wire \top/processor/sha_core/n340_135 ;
wire \top/processor/sha_core/n340_136 ;
wire \top/processor/sha_core/n340_137 ;
wire \top/processor/sha_core/n340_138 ;
wire \top/processor/sha_core/n340_139 ;
wire \top/processor/sha_core/n340_140 ;
wire \top/processor/sha_core/n340_141 ;
wire \top/processor/sha_core/n340_142 ;
wire \top/processor/sha_core/n340_143 ;
wire \top/processor/sha_core/n340_144 ;
wire \top/processor/sha_core/n340_145 ;
wire \top/processor/sha_core/n340_146 ;
wire \top/processor/sha_core/n340_147 ;
wire \top/processor/sha_core/n340_148 ;
wire \top/processor/sha_core/n340_149 ;
wire \top/processor/sha_core/n340_150 ;
wire \top/processor/sha_core/n340_151 ;
wire \top/processor/sha_core/n340_152 ;
wire \top/processor/sha_core/n340_153 ;
wire \top/processor/sha_core/n340_154 ;
wire \top/processor/sha_core/n340_155 ;
wire \top/processor/sha_core/n340_156 ;
wire \top/processor/sha_core/n340_157 ;
wire \top/processor/sha_core/n340_158 ;
wire \top/processor/sha_core/n340_159 ;
wire \top/processor/sha_core/n340_160 ;
wire \top/processor/sha_core/n340_161 ;
wire \top/processor/sha_core/n340_162 ;
wire \top/processor/sha_core/n340_163 ;
wire \top/processor/sha_core/n341_132 ;
wire \top/processor/sha_core/n341_133 ;
wire \top/processor/sha_core/n341_134 ;
wire \top/processor/sha_core/n341_135 ;
wire \top/processor/sha_core/n341_136 ;
wire \top/processor/sha_core/n341_137 ;
wire \top/processor/sha_core/n341_138 ;
wire \top/processor/sha_core/n341_139 ;
wire \top/processor/sha_core/n341_140 ;
wire \top/processor/sha_core/n341_141 ;
wire \top/processor/sha_core/n341_142 ;
wire \top/processor/sha_core/n341_143 ;
wire \top/processor/sha_core/n341_144 ;
wire \top/processor/sha_core/n341_145 ;
wire \top/processor/sha_core/n341_146 ;
wire \top/processor/sha_core/n341_147 ;
wire \top/processor/sha_core/n341_148 ;
wire \top/processor/sha_core/n341_149 ;
wire \top/processor/sha_core/n341_150 ;
wire \top/processor/sha_core/n341_151 ;
wire \top/processor/sha_core/n341_152 ;
wire \top/processor/sha_core/n341_153 ;
wire \top/processor/sha_core/n341_154 ;
wire \top/processor/sha_core/n341_155 ;
wire \top/processor/sha_core/n341_156 ;
wire \top/processor/sha_core/n341_157 ;
wire \top/processor/sha_core/n341_158 ;
wire \top/processor/sha_core/n341_159 ;
wire \top/processor/sha_core/n341_160 ;
wire \top/processor/sha_core/n341_161 ;
wire \top/processor/sha_core/n341_162 ;
wire \top/processor/sha_core/n341_163 ;
wire \top/processor/sha_core/n342_132 ;
wire \top/processor/sha_core/n342_133 ;
wire \top/processor/sha_core/n342_134 ;
wire \top/processor/sha_core/n342_135 ;
wire \top/processor/sha_core/n342_136 ;
wire \top/processor/sha_core/n342_137 ;
wire \top/processor/sha_core/n342_138 ;
wire \top/processor/sha_core/n342_139 ;
wire \top/processor/sha_core/n342_140 ;
wire \top/processor/sha_core/n342_141 ;
wire \top/processor/sha_core/n342_142 ;
wire \top/processor/sha_core/n342_143 ;
wire \top/processor/sha_core/n342_144 ;
wire \top/processor/sha_core/n342_145 ;
wire \top/processor/sha_core/n342_146 ;
wire \top/processor/sha_core/n342_147 ;
wire \top/processor/sha_core/n342_148 ;
wire \top/processor/sha_core/n342_149 ;
wire \top/processor/sha_core/n342_150 ;
wire \top/processor/sha_core/n342_151 ;
wire \top/processor/sha_core/n342_152 ;
wire \top/processor/sha_core/n342_153 ;
wire \top/processor/sha_core/n342_154 ;
wire \top/processor/sha_core/n342_155 ;
wire \top/processor/sha_core/n342_156 ;
wire \top/processor/sha_core/n342_157 ;
wire \top/processor/sha_core/n342_158 ;
wire \top/processor/sha_core/n342_159 ;
wire \top/processor/sha_core/n342_160 ;
wire \top/processor/sha_core/n342_161 ;
wire \top/processor/sha_core/n342_162 ;
wire \top/processor/sha_core/n342_163 ;
wire \top/processor/sha_core/n343_132 ;
wire \top/processor/sha_core/n343_133 ;
wire \top/processor/sha_core/n343_134 ;
wire \top/processor/sha_core/n343_135 ;
wire \top/processor/sha_core/n343_136 ;
wire \top/processor/sha_core/n343_137 ;
wire \top/processor/sha_core/n343_138 ;
wire \top/processor/sha_core/n343_139 ;
wire \top/processor/sha_core/n343_140 ;
wire \top/processor/sha_core/n343_141 ;
wire \top/processor/sha_core/n343_142 ;
wire \top/processor/sha_core/n343_143 ;
wire \top/processor/sha_core/n343_144 ;
wire \top/processor/sha_core/n343_145 ;
wire \top/processor/sha_core/n343_146 ;
wire \top/processor/sha_core/n343_147 ;
wire \top/processor/sha_core/n343_148 ;
wire \top/processor/sha_core/n343_149 ;
wire \top/processor/sha_core/n343_150 ;
wire \top/processor/sha_core/n343_151 ;
wire \top/processor/sha_core/n343_152 ;
wire \top/processor/sha_core/n343_153 ;
wire \top/processor/sha_core/n343_154 ;
wire \top/processor/sha_core/n343_155 ;
wire \top/processor/sha_core/n343_156 ;
wire \top/processor/sha_core/n343_157 ;
wire \top/processor/sha_core/n343_158 ;
wire \top/processor/sha_core/n343_159 ;
wire \top/processor/sha_core/n343_160 ;
wire \top/processor/sha_core/n343_161 ;
wire \top/processor/sha_core/n343_162 ;
wire \top/processor/sha_core/n343_163 ;
wire \top/processor/sha_core/n344_132 ;
wire \top/processor/sha_core/n344_133 ;
wire \top/processor/sha_core/n344_134 ;
wire \top/processor/sha_core/n344_135 ;
wire \top/processor/sha_core/n344_136 ;
wire \top/processor/sha_core/n344_137 ;
wire \top/processor/sha_core/n344_138 ;
wire \top/processor/sha_core/n344_139 ;
wire \top/processor/sha_core/n344_140 ;
wire \top/processor/sha_core/n344_141 ;
wire \top/processor/sha_core/n344_142 ;
wire \top/processor/sha_core/n344_143 ;
wire \top/processor/sha_core/n344_144 ;
wire \top/processor/sha_core/n344_145 ;
wire \top/processor/sha_core/n344_146 ;
wire \top/processor/sha_core/n344_147 ;
wire \top/processor/sha_core/n344_148 ;
wire \top/processor/sha_core/n344_149 ;
wire \top/processor/sha_core/n344_150 ;
wire \top/processor/sha_core/n344_151 ;
wire \top/processor/sha_core/n344_152 ;
wire \top/processor/sha_core/n344_153 ;
wire \top/processor/sha_core/n344_154 ;
wire \top/processor/sha_core/n344_155 ;
wire \top/processor/sha_core/n344_156 ;
wire \top/processor/sha_core/n344_157 ;
wire \top/processor/sha_core/n344_158 ;
wire \top/processor/sha_core/n344_159 ;
wire \top/processor/sha_core/n344_160 ;
wire \top/processor/sha_core/n344_161 ;
wire \top/processor/sha_core/n344_162 ;
wire \top/processor/sha_core/n344_163 ;
wire \top/processor/sha_core/n345_132 ;
wire \top/processor/sha_core/n345_133 ;
wire \top/processor/sha_core/n345_134 ;
wire \top/processor/sha_core/n345_135 ;
wire \top/processor/sha_core/n345_136 ;
wire \top/processor/sha_core/n345_137 ;
wire \top/processor/sha_core/n345_138 ;
wire \top/processor/sha_core/n345_139 ;
wire \top/processor/sha_core/n345_140 ;
wire \top/processor/sha_core/n345_141 ;
wire \top/processor/sha_core/n345_142 ;
wire \top/processor/sha_core/n345_143 ;
wire \top/processor/sha_core/n345_144 ;
wire \top/processor/sha_core/n345_145 ;
wire \top/processor/sha_core/n345_146 ;
wire \top/processor/sha_core/n345_147 ;
wire \top/processor/sha_core/n345_148 ;
wire \top/processor/sha_core/n345_149 ;
wire \top/processor/sha_core/n345_150 ;
wire \top/processor/sha_core/n345_151 ;
wire \top/processor/sha_core/n345_152 ;
wire \top/processor/sha_core/n345_153 ;
wire \top/processor/sha_core/n345_154 ;
wire \top/processor/sha_core/n345_155 ;
wire \top/processor/sha_core/n345_156 ;
wire \top/processor/sha_core/n345_157 ;
wire \top/processor/sha_core/n345_158 ;
wire \top/processor/sha_core/n345_159 ;
wire \top/processor/sha_core/n345_160 ;
wire \top/processor/sha_core/n345_161 ;
wire \top/processor/sha_core/n345_162 ;
wire \top/processor/sha_core/n345_163 ;
wire \top/processor/sha_core/n346_132 ;
wire \top/processor/sha_core/n346_133 ;
wire \top/processor/sha_core/n346_134 ;
wire \top/processor/sha_core/n346_135 ;
wire \top/processor/sha_core/n346_136 ;
wire \top/processor/sha_core/n346_137 ;
wire \top/processor/sha_core/n346_138 ;
wire \top/processor/sha_core/n346_139 ;
wire \top/processor/sha_core/n346_140 ;
wire \top/processor/sha_core/n346_141 ;
wire \top/processor/sha_core/n346_142 ;
wire \top/processor/sha_core/n346_143 ;
wire \top/processor/sha_core/n346_144 ;
wire \top/processor/sha_core/n346_145 ;
wire \top/processor/sha_core/n346_146 ;
wire \top/processor/sha_core/n346_147 ;
wire \top/processor/sha_core/n346_148 ;
wire \top/processor/sha_core/n346_149 ;
wire \top/processor/sha_core/n346_150 ;
wire \top/processor/sha_core/n346_151 ;
wire \top/processor/sha_core/n346_152 ;
wire \top/processor/sha_core/n346_153 ;
wire \top/processor/sha_core/n346_154 ;
wire \top/processor/sha_core/n346_155 ;
wire \top/processor/sha_core/n346_156 ;
wire \top/processor/sha_core/n346_157 ;
wire \top/processor/sha_core/n346_158 ;
wire \top/processor/sha_core/n346_159 ;
wire \top/processor/sha_core/n346_160 ;
wire \top/processor/sha_core/n346_161 ;
wire \top/processor/sha_core/n346_162 ;
wire \top/processor/sha_core/n346_163 ;
wire \top/processor/sha_core/n347_132 ;
wire \top/processor/sha_core/n347_133 ;
wire \top/processor/sha_core/n347_134 ;
wire \top/processor/sha_core/n347_135 ;
wire \top/processor/sha_core/n347_136 ;
wire \top/processor/sha_core/n347_137 ;
wire \top/processor/sha_core/n347_138 ;
wire \top/processor/sha_core/n347_139 ;
wire \top/processor/sha_core/n347_140 ;
wire \top/processor/sha_core/n347_141 ;
wire \top/processor/sha_core/n347_142 ;
wire \top/processor/sha_core/n347_143 ;
wire \top/processor/sha_core/n347_144 ;
wire \top/processor/sha_core/n347_145 ;
wire \top/processor/sha_core/n347_146 ;
wire \top/processor/sha_core/n347_147 ;
wire \top/processor/sha_core/n347_148 ;
wire \top/processor/sha_core/n347_149 ;
wire \top/processor/sha_core/n347_150 ;
wire \top/processor/sha_core/n347_151 ;
wire \top/processor/sha_core/n347_152 ;
wire \top/processor/sha_core/n347_153 ;
wire \top/processor/sha_core/n347_154 ;
wire \top/processor/sha_core/n347_155 ;
wire \top/processor/sha_core/n347_156 ;
wire \top/processor/sha_core/n347_157 ;
wire \top/processor/sha_core/n347_158 ;
wire \top/processor/sha_core/n347_159 ;
wire \top/processor/sha_core/n347_160 ;
wire \top/processor/sha_core/n347_161 ;
wire \top/processor/sha_core/n347_162 ;
wire \top/processor/sha_core/n347_163 ;
wire \top/processor/sha_core/n348_132 ;
wire \top/processor/sha_core/n348_133 ;
wire \top/processor/sha_core/n348_134 ;
wire \top/processor/sha_core/n348_135 ;
wire \top/processor/sha_core/n348_136 ;
wire \top/processor/sha_core/n348_137 ;
wire \top/processor/sha_core/n348_138 ;
wire \top/processor/sha_core/n348_139 ;
wire \top/processor/sha_core/n348_140 ;
wire \top/processor/sha_core/n348_141 ;
wire \top/processor/sha_core/n348_142 ;
wire \top/processor/sha_core/n348_143 ;
wire \top/processor/sha_core/n348_144 ;
wire \top/processor/sha_core/n348_145 ;
wire \top/processor/sha_core/n348_146 ;
wire \top/processor/sha_core/n348_147 ;
wire \top/processor/sha_core/n348_148 ;
wire \top/processor/sha_core/n348_149 ;
wire \top/processor/sha_core/n348_150 ;
wire \top/processor/sha_core/n348_151 ;
wire \top/processor/sha_core/n348_152 ;
wire \top/processor/sha_core/n348_153 ;
wire \top/processor/sha_core/n348_154 ;
wire \top/processor/sha_core/n348_155 ;
wire \top/processor/sha_core/n348_156 ;
wire \top/processor/sha_core/n348_157 ;
wire \top/processor/sha_core/n348_158 ;
wire \top/processor/sha_core/n348_159 ;
wire \top/processor/sha_core/n348_160 ;
wire \top/processor/sha_core/n348_161 ;
wire \top/processor/sha_core/n348_162 ;
wire \top/processor/sha_core/n348_163 ;
wire \top/processor/sha_core/n349_132 ;
wire \top/processor/sha_core/n349_133 ;
wire \top/processor/sha_core/n349_134 ;
wire \top/processor/sha_core/n349_135 ;
wire \top/processor/sha_core/n349_136 ;
wire \top/processor/sha_core/n349_137 ;
wire \top/processor/sha_core/n349_138 ;
wire \top/processor/sha_core/n349_139 ;
wire \top/processor/sha_core/n349_140 ;
wire \top/processor/sha_core/n349_141 ;
wire \top/processor/sha_core/n349_142 ;
wire \top/processor/sha_core/n349_143 ;
wire \top/processor/sha_core/n349_144 ;
wire \top/processor/sha_core/n349_145 ;
wire \top/processor/sha_core/n349_146 ;
wire \top/processor/sha_core/n349_147 ;
wire \top/processor/sha_core/n349_148 ;
wire \top/processor/sha_core/n349_149 ;
wire \top/processor/sha_core/n349_150 ;
wire \top/processor/sha_core/n349_151 ;
wire \top/processor/sha_core/n349_152 ;
wire \top/processor/sha_core/n349_153 ;
wire \top/processor/sha_core/n349_154 ;
wire \top/processor/sha_core/n349_155 ;
wire \top/processor/sha_core/n349_156 ;
wire \top/processor/sha_core/n349_157 ;
wire \top/processor/sha_core/n349_158 ;
wire \top/processor/sha_core/n349_159 ;
wire \top/processor/sha_core/n349_160 ;
wire \top/processor/sha_core/n349_161 ;
wire \top/processor/sha_core/n349_162 ;
wire \top/processor/sha_core/n349_163 ;
wire \top/processor/sha_core/n350_132 ;
wire \top/processor/sha_core/n350_133 ;
wire \top/processor/sha_core/n350_134 ;
wire \top/processor/sha_core/n350_135 ;
wire \top/processor/sha_core/n350_136 ;
wire \top/processor/sha_core/n350_137 ;
wire \top/processor/sha_core/n350_138 ;
wire \top/processor/sha_core/n350_139 ;
wire \top/processor/sha_core/n350_140 ;
wire \top/processor/sha_core/n350_141 ;
wire \top/processor/sha_core/n350_142 ;
wire \top/processor/sha_core/n350_143 ;
wire \top/processor/sha_core/n350_144 ;
wire \top/processor/sha_core/n350_145 ;
wire \top/processor/sha_core/n350_146 ;
wire \top/processor/sha_core/n350_147 ;
wire \top/processor/sha_core/n350_148 ;
wire \top/processor/sha_core/n350_149 ;
wire \top/processor/sha_core/n350_150 ;
wire \top/processor/sha_core/n350_151 ;
wire \top/processor/sha_core/n350_152 ;
wire \top/processor/sha_core/n350_153 ;
wire \top/processor/sha_core/n350_154 ;
wire \top/processor/sha_core/n350_155 ;
wire \top/processor/sha_core/n350_156 ;
wire \top/processor/sha_core/n350_157 ;
wire \top/processor/sha_core/n350_158 ;
wire \top/processor/sha_core/n350_159 ;
wire \top/processor/sha_core/n350_160 ;
wire \top/processor/sha_core/n350_161 ;
wire \top/processor/sha_core/n350_162 ;
wire \top/processor/sha_core/n350_163 ;
wire \top/processor/sha_core/n351_132 ;
wire \top/processor/sha_core/n351_133 ;
wire \top/processor/sha_core/n351_134 ;
wire \top/processor/sha_core/n351_135 ;
wire \top/processor/sha_core/n351_136 ;
wire \top/processor/sha_core/n351_137 ;
wire \top/processor/sha_core/n351_138 ;
wire \top/processor/sha_core/n351_139 ;
wire \top/processor/sha_core/n351_140 ;
wire \top/processor/sha_core/n351_141 ;
wire \top/processor/sha_core/n351_142 ;
wire \top/processor/sha_core/n351_143 ;
wire \top/processor/sha_core/n351_144 ;
wire \top/processor/sha_core/n351_145 ;
wire \top/processor/sha_core/n351_146 ;
wire \top/processor/sha_core/n351_147 ;
wire \top/processor/sha_core/n351_148 ;
wire \top/processor/sha_core/n351_149 ;
wire \top/processor/sha_core/n351_150 ;
wire \top/processor/sha_core/n351_151 ;
wire \top/processor/sha_core/n351_152 ;
wire \top/processor/sha_core/n351_153 ;
wire \top/processor/sha_core/n351_154 ;
wire \top/processor/sha_core/n351_155 ;
wire \top/processor/sha_core/n351_156 ;
wire \top/processor/sha_core/n351_157 ;
wire \top/processor/sha_core/n351_158 ;
wire \top/processor/sha_core/n351_159 ;
wire \top/processor/sha_core/n351_160 ;
wire \top/processor/sha_core/n351_161 ;
wire \top/processor/sha_core/n351_162 ;
wire \top/processor/sha_core/n351_163 ;
wire \top/processor/sha_core/n352_132 ;
wire \top/processor/sha_core/n352_133 ;
wire \top/processor/sha_core/n352_134 ;
wire \top/processor/sha_core/n352_135 ;
wire \top/processor/sha_core/n352_136 ;
wire \top/processor/sha_core/n352_137 ;
wire \top/processor/sha_core/n352_138 ;
wire \top/processor/sha_core/n352_139 ;
wire \top/processor/sha_core/n352_140 ;
wire \top/processor/sha_core/n352_141 ;
wire \top/processor/sha_core/n352_142 ;
wire \top/processor/sha_core/n352_143 ;
wire \top/processor/sha_core/n352_144 ;
wire \top/processor/sha_core/n352_145 ;
wire \top/processor/sha_core/n352_146 ;
wire \top/processor/sha_core/n352_147 ;
wire \top/processor/sha_core/n352_148 ;
wire \top/processor/sha_core/n352_149 ;
wire \top/processor/sha_core/n352_150 ;
wire \top/processor/sha_core/n352_151 ;
wire \top/processor/sha_core/n352_152 ;
wire \top/processor/sha_core/n352_153 ;
wire \top/processor/sha_core/n352_154 ;
wire \top/processor/sha_core/n352_155 ;
wire \top/processor/sha_core/n352_156 ;
wire \top/processor/sha_core/n352_157 ;
wire \top/processor/sha_core/n352_158 ;
wire \top/processor/sha_core/n352_159 ;
wire \top/processor/sha_core/n352_160 ;
wire \top/processor/sha_core/n352_161 ;
wire \top/processor/sha_core/n352_162 ;
wire \top/processor/sha_core/n352_163 ;
wire \top/processor/sha_core/n353_132 ;
wire \top/processor/sha_core/n353_133 ;
wire \top/processor/sha_core/n353_134 ;
wire \top/processor/sha_core/n353_135 ;
wire \top/processor/sha_core/n353_136 ;
wire \top/processor/sha_core/n353_137 ;
wire \top/processor/sha_core/n353_138 ;
wire \top/processor/sha_core/n353_139 ;
wire \top/processor/sha_core/n353_140 ;
wire \top/processor/sha_core/n353_141 ;
wire \top/processor/sha_core/n353_142 ;
wire \top/processor/sha_core/n353_143 ;
wire \top/processor/sha_core/n353_144 ;
wire \top/processor/sha_core/n353_145 ;
wire \top/processor/sha_core/n353_146 ;
wire \top/processor/sha_core/n353_147 ;
wire \top/processor/sha_core/n353_148 ;
wire \top/processor/sha_core/n353_149 ;
wire \top/processor/sha_core/n353_150 ;
wire \top/processor/sha_core/n353_151 ;
wire \top/processor/sha_core/n353_152 ;
wire \top/processor/sha_core/n353_153 ;
wire \top/processor/sha_core/n353_154 ;
wire \top/processor/sha_core/n353_155 ;
wire \top/processor/sha_core/n353_156 ;
wire \top/processor/sha_core/n353_157 ;
wire \top/processor/sha_core/n353_158 ;
wire \top/processor/sha_core/n353_159 ;
wire \top/processor/sha_core/n353_160 ;
wire \top/processor/sha_core/n353_161 ;
wire \top/processor/sha_core/n353_162 ;
wire \top/processor/sha_core/n353_163 ;
wire \top/processor/sha_core/n354_132 ;
wire \top/processor/sha_core/n354_133 ;
wire \top/processor/sha_core/n354_134 ;
wire \top/processor/sha_core/n354_135 ;
wire \top/processor/sha_core/n354_136 ;
wire \top/processor/sha_core/n354_137 ;
wire \top/processor/sha_core/n354_138 ;
wire \top/processor/sha_core/n354_139 ;
wire \top/processor/sha_core/n354_140 ;
wire \top/processor/sha_core/n354_141 ;
wire \top/processor/sha_core/n354_142 ;
wire \top/processor/sha_core/n354_143 ;
wire \top/processor/sha_core/n354_144 ;
wire \top/processor/sha_core/n354_145 ;
wire \top/processor/sha_core/n354_146 ;
wire \top/processor/sha_core/n354_147 ;
wire \top/processor/sha_core/n354_148 ;
wire \top/processor/sha_core/n354_149 ;
wire \top/processor/sha_core/n354_150 ;
wire \top/processor/sha_core/n354_151 ;
wire \top/processor/sha_core/n354_152 ;
wire \top/processor/sha_core/n354_153 ;
wire \top/processor/sha_core/n354_154 ;
wire \top/processor/sha_core/n354_155 ;
wire \top/processor/sha_core/n354_156 ;
wire \top/processor/sha_core/n354_157 ;
wire \top/processor/sha_core/n354_158 ;
wire \top/processor/sha_core/n354_159 ;
wire \top/processor/sha_core/n354_160 ;
wire \top/processor/sha_core/n354_161 ;
wire \top/processor/sha_core/n354_162 ;
wire \top/processor/sha_core/n354_163 ;
wire \top/processor/sha_core/n355_132 ;
wire \top/processor/sha_core/n355_133 ;
wire \top/processor/sha_core/n355_134 ;
wire \top/processor/sha_core/n355_135 ;
wire \top/processor/sha_core/n355_136 ;
wire \top/processor/sha_core/n355_137 ;
wire \top/processor/sha_core/n355_138 ;
wire \top/processor/sha_core/n355_139 ;
wire \top/processor/sha_core/n355_140 ;
wire \top/processor/sha_core/n355_141 ;
wire \top/processor/sha_core/n355_142 ;
wire \top/processor/sha_core/n355_143 ;
wire \top/processor/sha_core/n355_144 ;
wire \top/processor/sha_core/n355_145 ;
wire \top/processor/sha_core/n355_146 ;
wire \top/processor/sha_core/n355_147 ;
wire \top/processor/sha_core/n355_148 ;
wire \top/processor/sha_core/n355_149 ;
wire \top/processor/sha_core/n355_150 ;
wire \top/processor/sha_core/n355_151 ;
wire \top/processor/sha_core/n355_152 ;
wire \top/processor/sha_core/n355_153 ;
wire \top/processor/sha_core/n355_154 ;
wire \top/processor/sha_core/n355_155 ;
wire \top/processor/sha_core/n355_156 ;
wire \top/processor/sha_core/n355_157 ;
wire \top/processor/sha_core/n355_158 ;
wire \top/processor/sha_core/n355_159 ;
wire \top/processor/sha_core/n355_160 ;
wire \top/processor/sha_core/n355_161 ;
wire \top/processor/sha_core/n355_162 ;
wire \top/processor/sha_core/n355_163 ;
wire \top/processor/sha_core/n356_132 ;
wire \top/processor/sha_core/n356_133 ;
wire \top/processor/sha_core/n356_134 ;
wire \top/processor/sha_core/n356_135 ;
wire \top/processor/sha_core/n356_136 ;
wire \top/processor/sha_core/n356_137 ;
wire \top/processor/sha_core/n356_138 ;
wire \top/processor/sha_core/n356_139 ;
wire \top/processor/sha_core/n356_140 ;
wire \top/processor/sha_core/n356_141 ;
wire \top/processor/sha_core/n356_142 ;
wire \top/processor/sha_core/n356_143 ;
wire \top/processor/sha_core/n356_144 ;
wire \top/processor/sha_core/n356_145 ;
wire \top/processor/sha_core/n356_146 ;
wire \top/processor/sha_core/n356_147 ;
wire \top/processor/sha_core/n356_148 ;
wire \top/processor/sha_core/n356_149 ;
wire \top/processor/sha_core/n356_150 ;
wire \top/processor/sha_core/n356_151 ;
wire \top/processor/sha_core/n356_152 ;
wire \top/processor/sha_core/n356_153 ;
wire \top/processor/sha_core/n356_154 ;
wire \top/processor/sha_core/n356_155 ;
wire \top/processor/sha_core/n356_156 ;
wire \top/processor/sha_core/n356_157 ;
wire \top/processor/sha_core/n356_158 ;
wire \top/processor/sha_core/n356_159 ;
wire \top/processor/sha_core/n356_160 ;
wire \top/processor/sha_core/n356_161 ;
wire \top/processor/sha_core/n356_162 ;
wire \top/processor/sha_core/n356_163 ;
wire \top/processor/sha_core/n357_132 ;
wire \top/processor/sha_core/n357_133 ;
wire \top/processor/sha_core/n357_134 ;
wire \top/processor/sha_core/n357_135 ;
wire \top/processor/sha_core/n357_136 ;
wire \top/processor/sha_core/n357_137 ;
wire \top/processor/sha_core/n357_138 ;
wire \top/processor/sha_core/n357_139 ;
wire \top/processor/sha_core/n357_140 ;
wire \top/processor/sha_core/n357_141 ;
wire \top/processor/sha_core/n357_142 ;
wire \top/processor/sha_core/n357_143 ;
wire \top/processor/sha_core/n357_144 ;
wire \top/processor/sha_core/n357_145 ;
wire \top/processor/sha_core/n357_146 ;
wire \top/processor/sha_core/n357_147 ;
wire \top/processor/sha_core/n357_148 ;
wire \top/processor/sha_core/n357_149 ;
wire \top/processor/sha_core/n357_150 ;
wire \top/processor/sha_core/n357_151 ;
wire \top/processor/sha_core/n357_152 ;
wire \top/processor/sha_core/n357_153 ;
wire \top/processor/sha_core/n357_154 ;
wire \top/processor/sha_core/n357_155 ;
wire \top/processor/sha_core/n357_156 ;
wire \top/processor/sha_core/n357_157 ;
wire \top/processor/sha_core/n357_158 ;
wire \top/processor/sha_core/n357_159 ;
wire \top/processor/sha_core/n357_160 ;
wire \top/processor/sha_core/n357_161 ;
wire \top/processor/sha_core/n357_162 ;
wire \top/processor/sha_core/n357_163 ;
wire \top/processor/sha_core/n358_132 ;
wire \top/processor/sha_core/n358_133 ;
wire \top/processor/sha_core/n358_134 ;
wire \top/processor/sha_core/n358_135 ;
wire \top/processor/sha_core/n358_136 ;
wire \top/processor/sha_core/n358_137 ;
wire \top/processor/sha_core/n358_138 ;
wire \top/processor/sha_core/n358_139 ;
wire \top/processor/sha_core/n358_140 ;
wire \top/processor/sha_core/n358_141 ;
wire \top/processor/sha_core/n358_142 ;
wire \top/processor/sha_core/n358_143 ;
wire \top/processor/sha_core/n358_144 ;
wire \top/processor/sha_core/n358_145 ;
wire \top/processor/sha_core/n358_146 ;
wire \top/processor/sha_core/n358_147 ;
wire \top/processor/sha_core/n358_148 ;
wire \top/processor/sha_core/n358_149 ;
wire \top/processor/sha_core/n358_150 ;
wire \top/processor/sha_core/n358_151 ;
wire \top/processor/sha_core/n358_152 ;
wire \top/processor/sha_core/n358_153 ;
wire \top/processor/sha_core/n358_154 ;
wire \top/processor/sha_core/n358_155 ;
wire \top/processor/sha_core/n358_156 ;
wire \top/processor/sha_core/n358_157 ;
wire \top/processor/sha_core/n358_158 ;
wire \top/processor/sha_core/n358_159 ;
wire \top/processor/sha_core/n358_160 ;
wire \top/processor/sha_core/n358_161 ;
wire \top/processor/sha_core/n358_162 ;
wire \top/processor/sha_core/n358_163 ;
wire \top/processor/sha_core/n36_3 ;
wire \top/processor/sha_core/n37_3 ;
wire \top/processor/sha_core/n38_3 ;
wire \top/processor/sha_core/n39_3 ;
wire \top/processor/sha_core/n40_3 ;
wire \top/processor/sha_core/n41_3 ;
wire \top/processor/sha_core/n42_3 ;
wire \top/processor/sha_core/n43_3 ;
wire \top/processor/sha_core/n44_3 ;
wire \top/processor/sha_core/n45_3 ;
wire \top/processor/sha_core/n46_3 ;
wire \top/processor/sha_core/n47_3 ;
wire \top/processor/sha_core/n48_3 ;
wire \top/processor/sha_core/n49_3 ;
wire \top/processor/sha_core/n50_3 ;
wire \top/processor/sha_core/n51_3 ;
wire \top/processor/sha_core/n52_3 ;
wire \top/processor/sha_core/n53_3 ;
wire \top/processor/sha_core/n54_3 ;
wire \top/processor/sha_core/n55_3 ;
wire \top/processor/sha_core/n56_3 ;
wire \top/processor/sha_core/n57_3 ;
wire \top/processor/sha_core/n58_3 ;
wire \top/processor/sha_core/n59_3 ;
wire \top/processor/sha_core/n60_3 ;
wire \top/processor/sha_core/n61_3 ;
wire \top/processor/sha_core/n62_3 ;
wire \top/processor/sha_core/n63_3 ;
wire \top/processor/sha_core/n64_3 ;
wire \top/processor/sha_core/n65_3 ;
wire \top/processor/sha_core/n66_3 ;
wire \top/processor/sha_core/n67_3 ;
wire \top/processor/sha_core/n197_3 ;
wire \top/processor/sha_core/n198_3 ;
wire \top/processor/sha_core/n199_3 ;
wire \top/processor/sha_core/n200_3 ;
wire \top/processor/sha_core/n201_3 ;
wire \top/processor/sha_core/n202_3 ;
wire \top/processor/sha_core/n203_3 ;
wire \top/processor/sha_core/n204_3 ;
wire \top/processor/sha_core/n205_3 ;
wire \top/processor/sha_core/n206_3 ;
wire \top/processor/sha_core/n207_3 ;
wire \top/processor/sha_core/n208_3 ;
wire \top/processor/sha_core/n209_3 ;
wire \top/processor/sha_core/n210_3 ;
wire \top/processor/sha_core/n211_3 ;
wire \top/processor/sha_core/n212_3 ;
wire \top/processor/sha_core/n213_3 ;
wire \top/processor/sha_core/n214_3 ;
wire \top/processor/sha_core/n215_3 ;
wire \top/processor/sha_core/n216_3 ;
wire \top/processor/sha_core/n217_3 ;
wire \top/processor/sha_core/n218_3 ;
wire \top/processor/sha_core/n219_3 ;
wire \top/processor/sha_core/n220_3 ;
wire \top/processor/sha_core/n221_3 ;
wire \top/processor/sha_core/n222_3 ;
wire \top/processor/sha_core/n223_3 ;
wire \top/processor/sha_core/n224_3 ;
wire \top/processor/sha_core/n225_3 ;
wire \top/processor/sha_core/n226_3 ;
wire \top/processor/sha_core/n227_3 ;
wire \top/processor/sha_core/n228_3 ;
wire \top/processor/sha_core/n424_3 ;
wire \top/processor/sha_core/n425_3 ;
wire \top/processor/sha_core/n426_3 ;
wire \top/processor/sha_core/n427_3 ;
wire \top/processor/sha_core/n428_3 ;
wire \top/processor/sha_core/n429_3 ;
wire \top/processor/sha_core/n430_3 ;
wire \top/processor/sha_core/n431_3 ;
wire \top/processor/sha_core/n432_3 ;
wire \top/processor/sha_core/n433_3 ;
wire \top/processor/sha_core/n434_3 ;
wire \top/processor/sha_core/n435_3 ;
wire \top/processor/sha_core/n436_3 ;
wire \top/processor/sha_core/n437_3 ;
wire \top/processor/sha_core/n438_3 ;
wire \top/processor/sha_core/n439_3 ;
wire \top/processor/sha_core/n440_3 ;
wire \top/processor/sha_core/n441_3 ;
wire \top/processor/sha_core/n442_3 ;
wire \top/processor/sha_core/n443_3 ;
wire \top/processor/sha_core/n444_3 ;
wire \top/processor/sha_core/n445_3 ;
wire \top/processor/sha_core/n446_3 ;
wire \top/processor/sha_core/n447_3 ;
wire \top/processor/sha_core/n448_3 ;
wire \top/processor/sha_core/n449_3 ;
wire \top/processor/sha_core/n450_3 ;
wire \top/processor/sha_core/n451_3 ;
wire \top/processor/sha_core/n452_3 ;
wire \top/processor/sha_core/n453_3 ;
wire \top/processor/sha_core/n454_3 ;
wire \top/processor/sha_core/n455_3 ;
wire \top/processor/sha_core/n584_3 ;
wire \top/processor/sha_core/n585_3 ;
wire \top/processor/sha_core/n586_3 ;
wire \top/processor/sha_core/n587_3 ;
wire \top/processor/sha_core/n588_3 ;
wire \top/processor/sha_core/n589_3 ;
wire \top/processor/sha_core/n590_3 ;
wire \top/processor/sha_core/n591_3 ;
wire \top/processor/sha_core/n592_3 ;
wire \top/processor/sha_core/n593_3 ;
wire \top/processor/sha_core/n594_3 ;
wire \top/processor/sha_core/n595_3 ;
wire \top/processor/sha_core/n596_3 ;
wire \top/processor/sha_core/n597_3 ;
wire \top/processor/sha_core/n598_3 ;
wire \top/processor/sha_core/n599_3 ;
wire \top/processor/sha_core/n600_3 ;
wire \top/processor/sha_core/n601_3 ;
wire \top/processor/sha_core/n602_3 ;
wire \top/processor/sha_core/n603_3 ;
wire \top/processor/sha_core/n604_3 ;
wire \top/processor/sha_core/n605_3 ;
wire \top/processor/sha_core/n606_3 ;
wire \top/processor/sha_core/n607_3 ;
wire \top/processor/sha_core/n608_3 ;
wire \top/processor/sha_core/n609_3 ;
wire \top/processor/sha_core/n610_3 ;
wire \top/processor/sha_core/n611_3 ;
wire \top/processor/sha_core/n612_3 ;
wire \top/processor/sha_core/n613_3 ;
wire \top/processor/sha_core/n614_3 ;
wire \top/processor/sha_core/n615_3 ;
wire \top/processor/sha_core/n3543_3 ;
wire \top/processor/sha_core/n3545_3 ;
wire \top/processor/sha_core/n3546_3 ;
wire \top/processor/sha_core/n3547_3 ;
wire \top/processor/sha_core/n3548_3 ;
wire \top/processor/sha_core/n3549_3 ;
wire \top/processor/sha_core/n3550_3 ;
wire \top/processor/sha_core/n3551_3 ;
wire \top/processor/sha_core/n3552_3 ;
wire \top/processor/sha_core/n3553_3 ;
wire \top/processor/sha_core/n3554_3 ;
wire \top/processor/sha_core/n3555_3 ;
wire \top/processor/sha_core/n3556_3 ;
wire \top/processor/sha_core/n3557_3 ;
wire \top/processor/sha_core/n3558_3 ;
wire \top/processor/sha_core/n3559_3 ;
wire \top/processor/sha_core/n3560_3 ;
wire \top/processor/sha_core/n3561_3 ;
wire \top/processor/sha_core/n3562_3 ;
wire \top/processor/sha_core/n3563_3 ;
wire \top/processor/sha_core/n3564_3 ;
wire \top/processor/sha_core/n3565_3 ;
wire \top/processor/sha_core/n3566_3 ;
wire \top/processor/sha_core/n3567_3 ;
wire \top/processor/sha_core/n3568_3 ;
wire \top/processor/sha_core/n3569_3 ;
wire \top/processor/sha_core/n3570_3 ;
wire \top/processor/sha_core/n3571_3 ;
wire \top/processor/sha_core/n3572_3 ;
wire \top/processor/sha_core/n3573_3 ;
wire \top/processor/sha_core/n3769_3 ;
wire \top/processor/sha_core/n3770_3 ;
wire \top/processor/sha_core/n3771_3 ;
wire \top/processor/sha_core/n3772_3 ;
wire \top/processor/sha_core/n3773_3 ;
wire \top/processor/sha_core/n3774_3 ;
wire \top/processor/sha_core/n3775_3 ;
wire \top/processor/sha_core/n3776_3 ;
wire \top/processor/sha_core/n3777_3 ;
wire \top/processor/sha_core/n3778_3 ;
wire \top/processor/sha_core/n3779_3 ;
wire \top/processor/sha_core/n3780_3 ;
wire \top/processor/sha_core/n3781_3 ;
wire \top/processor/sha_core/n3782_3 ;
wire \top/processor/sha_core/n3783_3 ;
wire \top/processor/sha_core/n3784_3 ;
wire \top/processor/sha_core/n3785_3 ;
wire \top/processor/sha_core/n3786_3 ;
wire \top/processor/sha_core/n3787_3 ;
wire \top/processor/sha_core/n3788_3 ;
wire \top/processor/sha_core/n3789_3 ;
wire \top/processor/sha_core/n3790_3 ;
wire \top/processor/sha_core/n3791_3 ;
wire \top/processor/sha_core/n3792_3 ;
wire \top/processor/sha_core/n3793_3 ;
wire \top/processor/sha_core/n3794_3 ;
wire \top/processor/sha_core/n3795_3 ;
wire \top/processor/sha_core/n3796_3 ;
wire \top/processor/sha_core/n3797_3 ;
wire \top/processor/sha_core/n8430_3 ;
wire \top/processor/sha_core/n8431_3 ;
wire \top/processor/sha_core/n8432_3 ;
wire \top/processor/sha_core/n8433_3 ;
wire \top/processor/sha_core/n8434_3 ;
wire \top/processor/sha_core/n8435_3 ;
wire \top/processor/sha_core/n8436_3 ;
wire \top/processor/sha_core/n8437_3 ;
wire \top/processor/sha_core/n8438_3 ;
wire \top/processor/sha_core/n8439_3 ;
wire \top/processor/sha_core/n8440_3 ;
wire \top/processor/sha_core/n8441_3 ;
wire \top/processor/sha_core/n8442_3 ;
wire \top/processor/sha_core/n8443_3 ;
wire \top/processor/sha_core/n8444_3 ;
wire \top/processor/sha_core/n8445_3 ;
wire \top/processor/sha_core/n8446_3 ;
wire \top/processor/sha_core/n8447_3 ;
wire \top/processor/sha_core/n8448_3 ;
wire \top/processor/sha_core/n8449_3 ;
wire \top/processor/sha_core/n8450_3 ;
wire \top/processor/sha_core/n8451_3 ;
wire \top/processor/sha_core/n8452_3 ;
wire \top/processor/sha_core/n8453_3 ;
wire \top/processor/sha_core/n8454_3 ;
wire \top/processor/sha_core/n8455_3 ;
wire \top/processor/sha_core/n8456_3 ;
wire \top/processor/sha_core/n8457_3 ;
wire \top/processor/sha_core/n8458_3 ;
wire \top/processor/sha_core/n8459_3 ;
wire \top/processor/sha_core/n8460_3 ;
wire \top/processor/sha_core/n8461_3 ;
wire \top/processor/sha_core/n11869_11 ;
wire \top/processor/sha_core/n11872_9 ;
wire \top/processor/sha_core/n11873_9 ;
wire \top/processor/sha_core/n11874_9 ;
wire \top/processor/sha_core/n11875_9 ;
wire \top/processor/sha_core/n11876_9 ;
wire \top/processor/sha_core/n11877_9 ;
wire \top/processor/sha_core/n11878_9 ;
wire \top/processor/sha_core/n11879_9 ;
wire \top/processor/sha_core/n11880_9 ;
wire \top/processor/sha_core/n11881_9 ;
wire \top/processor/sha_core/n11882_9 ;
wire \top/processor/sha_core/n11883_9 ;
wire \top/processor/sha_core/n11884_9 ;
wire \top/processor/sha_core/n11885_9 ;
wire \top/processor/sha_core/n11886_9 ;
wire \top/processor/sha_core/n11887_9 ;
wire \top/processor/sha_core/n11888_9 ;
wire \top/processor/sha_core/n11889_9 ;
wire \top/processor/sha_core/n11890_9 ;
wire \top/processor/sha_core/n11891_9 ;
wire \top/processor/sha_core/n11892_9 ;
wire \top/processor/sha_core/n11893_9 ;
wire \top/processor/sha_core/n11894_9 ;
wire \top/processor/sha_core/n11895_9 ;
wire \top/processor/sha_core/n11896_9 ;
wire \top/processor/sha_core/n11897_9 ;
wire \top/processor/sha_core/n11898_9 ;
wire \top/processor/sha_core/n11899_9 ;
wire \top/processor/sha_core/n11900_9 ;
wire \top/processor/sha_core/n11901_9 ;
wire \top/processor/sha_core/n11902_9 ;
wire \top/processor/sha_core/n11903_9 ;
wire \top/processor/sha_core/n11904_9 ;
wire \top/processor/sha_core/n11905_9 ;
wire \top/processor/sha_core/n11906_9 ;
wire \top/processor/sha_core/n11907_9 ;
wire \top/processor/sha_core/n11908_9 ;
wire \top/processor/sha_core/n11909_9 ;
wire \top/processor/sha_core/n11910_9 ;
wire \top/processor/sha_core/n11911_9 ;
wire \top/processor/sha_core/n11912_9 ;
wire \top/processor/sha_core/n11913_9 ;
wire \top/processor/sha_core/n11914_9 ;
wire \top/processor/sha_core/n11915_9 ;
wire \top/processor/sha_core/n11916_9 ;
wire \top/processor/sha_core/n11917_9 ;
wire \top/processor/sha_core/n11918_9 ;
wire \top/processor/sha_core/n11919_9 ;
wire \top/processor/sha_core/n11920_9 ;
wire \top/processor/sha_core/n11921_9 ;
wire \top/processor/sha_core/n11922_9 ;
wire \top/processor/sha_core/n11923_9 ;
wire \top/processor/sha_core/n11924_9 ;
wire \top/processor/sha_core/n11925_9 ;
wire \top/processor/sha_core/n11926_9 ;
wire \top/processor/sha_core/n11927_9 ;
wire \top/processor/sha_core/n11928_9 ;
wire \top/processor/sha_core/n11929_9 ;
wire \top/processor/sha_core/n11930_9 ;
wire \top/processor/sha_core/n11931_9 ;
wire \top/processor/sha_core/n11932_9 ;
wire \top/processor/sha_core/n11933_9 ;
wire \top/processor/sha_core/n11934_9 ;
wire \top/processor/sha_core/n11935_9 ;
wire \top/processor/sha_core/n11936_9 ;
wire \top/processor/sha_core/n11937_9 ;
wire \top/processor/sha_core/n11938_9 ;
wire \top/processor/sha_core/n11939_9 ;
wire \top/processor/sha_core/n11940_9 ;
wire \top/processor/sha_core/n11941_9 ;
wire \top/processor/sha_core/n11942_9 ;
wire \top/processor/sha_core/n11943_9 ;
wire \top/processor/sha_core/n11944_9 ;
wire \top/processor/sha_core/n11945_9 ;
wire \top/processor/sha_core/n11946_9 ;
wire \top/processor/sha_core/n11947_9 ;
wire \top/processor/sha_core/n11948_9 ;
wire \top/processor/sha_core/n11949_9 ;
wire \top/processor/sha_core/n11950_9 ;
wire \top/processor/sha_core/n11951_9 ;
wire \top/processor/sha_core/n11952_9 ;
wire \top/processor/sha_core/n11953_9 ;
wire \top/processor/sha_core/n11954_9 ;
wire \top/processor/sha_core/n11955_9 ;
wire \top/processor/sha_core/n11956_9 ;
wire \top/processor/sha_core/n11957_9 ;
wire \top/processor/sha_core/n11958_9 ;
wire \top/processor/sha_core/n11959_9 ;
wire \top/processor/sha_core/n11960_9 ;
wire \top/processor/sha_core/n11961_9 ;
wire \top/processor/sha_core/n11962_9 ;
wire \top/processor/sha_core/n11963_9 ;
wire \top/processor/sha_core/n11964_9 ;
wire \top/processor/sha_core/n11965_9 ;
wire \top/processor/sha_core/n11966_9 ;
wire \top/processor/sha_core/n11967_9 ;
wire \top/processor/sha_core/n11968_9 ;
wire \top/processor/sha_core/n11969_9 ;
wire \top/processor/sha_core/n11970_9 ;
wire \top/processor/sha_core/n11971_9 ;
wire \top/processor/sha_core/n11972_9 ;
wire \top/processor/sha_core/n11973_9 ;
wire \top/processor/sha_core/n11974_9 ;
wire \top/processor/sha_core/n11975_9 ;
wire \top/processor/sha_core/n11976_9 ;
wire \top/processor/sha_core/n11977_9 ;
wire \top/processor/sha_core/n11978_9 ;
wire \top/processor/sha_core/n11979_9 ;
wire \top/processor/sha_core/n11980_9 ;
wire \top/processor/sha_core/n11981_9 ;
wire \top/processor/sha_core/n11982_9 ;
wire \top/processor/sha_core/n11983_9 ;
wire \top/processor/sha_core/n11984_9 ;
wire \top/processor/sha_core/n11985_9 ;
wire \top/processor/sha_core/n11986_9 ;
wire \top/processor/sha_core/n11987_9 ;
wire \top/processor/sha_core/n11988_9 ;
wire \top/processor/sha_core/n11989_9 ;
wire \top/processor/sha_core/n11990_9 ;
wire \top/processor/sha_core/n11991_9 ;
wire \top/processor/sha_core/n11992_9 ;
wire \top/processor/sha_core/n11993_9 ;
wire \top/processor/sha_core/n11994_9 ;
wire \top/processor/sha_core/n11995_9 ;
wire \top/processor/sha_core/n11996_9 ;
wire \top/processor/sha_core/n11997_9 ;
wire \top/processor/sha_core/n11998_9 ;
wire \top/processor/sha_core/n11999_9 ;
wire \top/processor/sha_core/n12000_9 ;
wire \top/processor/sha_core/n12001_9 ;
wire \top/processor/sha_core/n12002_9 ;
wire \top/processor/sha_core/n12003_9 ;
wire \top/processor/sha_core/n12004_9 ;
wire \top/processor/sha_core/n12005_9 ;
wire \top/processor/sha_core/n12006_9 ;
wire \top/processor/sha_core/n12007_9 ;
wire \top/processor/sha_core/n12008_9 ;
wire \top/processor/sha_core/n12009_9 ;
wire \top/processor/sha_core/n12010_9 ;
wire \top/processor/sha_core/n12011_9 ;
wire \top/processor/sha_core/n12012_9 ;
wire \top/processor/sha_core/n12013_9 ;
wire \top/processor/sha_core/n12014_9 ;
wire \top/processor/sha_core/n12015_9 ;
wire \top/processor/sha_core/n12016_9 ;
wire \top/processor/sha_core/n12017_9 ;
wire \top/processor/sha_core/n12018_9 ;
wire \top/processor/sha_core/n12019_9 ;
wire \top/processor/sha_core/n12020_9 ;
wire \top/processor/sha_core/n12021_9 ;
wire \top/processor/sha_core/n12022_9 ;
wire \top/processor/sha_core/n12023_9 ;
wire \top/processor/sha_core/n12024_9 ;
wire \top/processor/sha_core/n12025_9 ;
wire \top/processor/sha_core/n12026_9 ;
wire \top/processor/sha_core/n12027_9 ;
wire \top/processor/sha_core/n12028_9 ;
wire \top/processor/sha_core/n12029_9 ;
wire \top/processor/sha_core/n12030_9 ;
wire \top/processor/sha_core/n12031_9 ;
wire \top/processor/sha_core/n12032_9 ;
wire \top/processor/sha_core/n12033_9 ;
wire \top/processor/sha_core/n12034_9 ;
wire \top/processor/sha_core/n12035_9 ;
wire \top/processor/sha_core/n12036_9 ;
wire \top/processor/sha_core/n12037_9 ;
wire \top/processor/sha_core/n12038_9 ;
wire \top/processor/sha_core/n12039_9 ;
wire \top/processor/sha_core/n12040_9 ;
wire \top/processor/sha_core/n12041_9 ;
wire \top/processor/sha_core/n12042_9 ;
wire \top/processor/sha_core/n12043_9 ;
wire \top/processor/sha_core/n12044_9 ;
wire \top/processor/sha_core/n12045_9 ;
wire \top/processor/sha_core/n12046_9 ;
wire \top/processor/sha_core/n12047_9 ;
wire \top/processor/sha_core/n12048_9 ;
wire \top/processor/sha_core/n12049_9 ;
wire \top/processor/sha_core/n12050_9 ;
wire \top/processor/sha_core/n12051_9 ;
wire \top/processor/sha_core/n12052_9 ;
wire \top/processor/sha_core/n12053_9 ;
wire \top/processor/sha_core/n12054_9 ;
wire \top/processor/sha_core/n12055_9 ;
wire \top/processor/sha_core/n12056_9 ;
wire \top/processor/sha_core/n12057_9 ;
wire \top/processor/sha_core/n12058_9 ;
wire \top/processor/sha_core/n12059_9 ;
wire \top/processor/sha_core/n12060_9 ;
wire \top/processor/sha_core/n12061_9 ;
wire \top/processor/sha_core/n12062_9 ;
wire \top/processor/sha_core/n12063_9 ;
wire \top/processor/sha_core/n12064_9 ;
wire \top/processor/sha_core/n12065_9 ;
wire \top/processor/sha_core/n12066_9 ;
wire \top/processor/sha_core/n12067_9 ;
wire \top/processor/sha_core/n12068_9 ;
wire \top/processor/sha_core/n12069_9 ;
wire \top/processor/sha_core/n12070_9 ;
wire \top/processor/sha_core/n12071_9 ;
wire \top/processor/sha_core/n12072_9 ;
wire \top/processor/sha_core/n12073_9 ;
wire \top/processor/sha_core/n12074_9 ;
wire \top/processor/sha_core/n12075_9 ;
wire \top/processor/sha_core/n12076_9 ;
wire \top/processor/sha_core/n12077_9 ;
wire \top/processor/sha_core/n12078_9 ;
wire \top/processor/sha_core/n12079_9 ;
wire \top/processor/sha_core/n12080_9 ;
wire \top/processor/sha_core/n12081_9 ;
wire \top/processor/sha_core/n12082_9 ;
wire \top/processor/sha_core/n12083_9 ;
wire \top/processor/sha_core/n12084_9 ;
wire \top/processor/sha_core/n12085_9 ;
wire \top/processor/sha_core/n12086_9 ;
wire \top/processor/sha_core/n12087_9 ;
wire \top/processor/sha_core/n12088_9 ;
wire \top/processor/sha_core/n12089_9 ;
wire \top/processor/sha_core/n12090_9 ;
wire \top/processor/sha_core/n12091_9 ;
wire \top/processor/sha_core/n12092_9 ;
wire \top/processor/sha_core/n12093_9 ;
wire \top/processor/sha_core/n12094_9 ;
wire \top/processor/sha_core/n12095_9 ;
wire \top/processor/sha_core/n12096_9 ;
wire \top/processor/sha_core/n12097_9 ;
wire \top/processor/sha_core/n12098_9 ;
wire \top/processor/sha_core/n12099_9 ;
wire \top/processor/sha_core/n12100_9 ;
wire \top/processor/sha_core/n12101_9 ;
wire \top/processor/sha_core/n12102_9 ;
wire \top/processor/sha_core/n12103_9 ;
wire \top/processor/sha_core/n12104_9 ;
wire \top/processor/sha_core/n12105_9 ;
wire \top/processor/sha_core/n12106_9 ;
wire \top/processor/sha_core/n12107_9 ;
wire \top/processor/sha_core/n12108_9 ;
wire \top/processor/sha_core/n12109_9 ;
wire \top/processor/sha_core/n12110_9 ;
wire \top/processor/sha_core/n12111_9 ;
wire \top/processor/sha_core/n12112_9 ;
wire \top/processor/sha_core/n12113_9 ;
wire \top/processor/sha_core/n12114_9 ;
wire \top/processor/sha_core/n12115_9 ;
wire \top/processor/sha_core/n12116_9 ;
wire \top/processor/sha_core/n12117_9 ;
wire \top/processor/sha_core/n12118_9 ;
wire \top/processor/sha_core/n12119_9 ;
wire \top/processor/sha_core/n12120_9 ;
wire \top/processor/sha_core/n12121_9 ;
wire \top/processor/sha_core/n12122_9 ;
wire \top/processor/sha_core/n12123_9 ;
wire \top/processor/sha_core/n12124_9 ;
wire \top/processor/sha_core/n12125_9 ;
wire \top/processor/sha_core/n12126_9 ;
wire \top/processor/sha_core/n12127_9 ;
wire \top/processor/sha_core/n12135_10 ;
wire \top/processor/sha_core/n12136_9 ;
wire \top/processor/sha_core/n12137_9 ;
wire \top/processor/sha_core/n12138_9 ;
wire \top/processor/sha_core/n12139_9 ;
wire \top/processor/sha_core/n12140_9 ;
wire \top/processor/sha_core/n12141_9 ;
wire \top/processor/sha_core/n12142_9 ;
wire \top/processor/sha_core/n12143_9 ;
wire \top/processor/sha_core/n12144_9 ;
wire \top/processor/sha_core/n12145_9 ;
wire \top/processor/sha_core/n12146_9 ;
wire \top/processor/sha_core/n12147_9 ;
wire \top/processor/sha_core/n12148_9 ;
wire \top/processor/sha_core/n12149_9 ;
wire \top/processor/sha_core/n12150_9 ;
wire \top/processor/sha_core/n12151_9 ;
wire \top/processor/sha_core/n12152_9 ;
wire \top/processor/sha_core/n12153_9 ;
wire \top/processor/sha_core/n12154_9 ;
wire \top/processor/sha_core/n12155_9 ;
wire \top/processor/sha_core/n12156_9 ;
wire \top/processor/sha_core/n12157_9 ;
wire \top/processor/sha_core/n12158_9 ;
wire \top/processor/sha_core/n12159_9 ;
wire \top/processor/sha_core/n12160_9 ;
wire \top/processor/sha_core/n12161_9 ;
wire \top/processor/sha_core/n12162_9 ;
wire \top/processor/sha_core/n12163_9 ;
wire \top/processor/sha_core/n12164_9 ;
wire \top/processor/sha_core/n12165_9 ;
wire \top/processor/sha_core/n12166_9 ;
wire \top/processor/sha_core/n12167_9 ;
wire \top/processor/sha_core/n12168_9 ;
wire \top/processor/sha_core/n12169_9 ;
wire \top/processor/sha_core/n12170_9 ;
wire \top/processor/sha_core/n12171_9 ;
wire \top/processor/sha_core/n12172_9 ;
wire \top/processor/sha_core/n12173_9 ;
wire \top/processor/sha_core/n12174_9 ;
wire \top/processor/sha_core/n12175_9 ;
wire \top/processor/sha_core/n12176_9 ;
wire \top/processor/sha_core/n12177_9 ;
wire \top/processor/sha_core/n12178_9 ;
wire \top/processor/sha_core/n12179_9 ;
wire \top/processor/sha_core/n12180_9 ;
wire \top/processor/sha_core/n12181_9 ;
wire \top/processor/sha_core/n12182_9 ;
wire \top/processor/sha_core/n12183_9 ;
wire \top/processor/sha_core/n12184_9 ;
wire \top/processor/sha_core/n12185_9 ;
wire \top/processor/sha_core/n12186_9 ;
wire \top/processor/sha_core/n12187_9 ;
wire \top/processor/sha_core/n12188_9 ;
wire \top/processor/sha_core/n12189_9 ;
wire \top/processor/sha_core/n12190_9 ;
wire \top/processor/sha_core/n12191_9 ;
wire \top/processor/sha_core/n12192_9 ;
wire \top/processor/sha_core/n12193_9 ;
wire \top/processor/sha_core/n12194_9 ;
wire \top/processor/sha_core/n12195_9 ;
wire \top/processor/sha_core/n12196_9 ;
wire \top/processor/sha_core/n12197_9 ;
wire \top/processor/sha_core/n12198_9 ;
wire \top/processor/sha_core/n12199_9 ;
wire \top/processor/sha_core/n12200_9 ;
wire \top/processor/sha_core/n12201_9 ;
wire \top/processor/sha_core/n12202_9 ;
wire \top/processor/sha_core/n12203_9 ;
wire \top/processor/sha_core/n12204_9 ;
wire \top/processor/sha_core/n12205_9 ;
wire \top/processor/sha_core/n12206_9 ;
wire \top/processor/sha_core/n12207_9 ;
wire \top/processor/sha_core/n12208_9 ;
wire \top/processor/sha_core/n12209_9 ;
wire \top/processor/sha_core/n12210_9 ;
wire \top/processor/sha_core/n12211_9 ;
wire \top/processor/sha_core/n12212_9 ;
wire \top/processor/sha_core/n12213_9 ;
wire \top/processor/sha_core/n12214_9 ;
wire \top/processor/sha_core/n12215_9 ;
wire \top/processor/sha_core/n12216_9 ;
wire \top/processor/sha_core/n12217_9 ;
wire \top/processor/sha_core/n12218_9 ;
wire \top/processor/sha_core/n12219_9 ;
wire \top/processor/sha_core/n12220_9 ;
wire \top/processor/sha_core/n12221_9 ;
wire \top/processor/sha_core/n12222_9 ;
wire \top/processor/sha_core/n12223_9 ;
wire \top/processor/sha_core/n12224_9 ;
wire \top/processor/sha_core/n12225_9 ;
wire \top/processor/sha_core/n12226_9 ;
wire \top/processor/sha_core/n12227_9 ;
wire \top/processor/sha_core/n12228_9 ;
wire \top/processor/sha_core/n12229_9 ;
wire \top/processor/sha_core/n12230_9 ;
wire \top/processor/sha_core/n12231_9 ;
wire \top/processor/sha_core/n12232_9 ;
wire \top/processor/sha_core/n12233_9 ;
wire \top/processor/sha_core/n12234_9 ;
wire \top/processor/sha_core/n12235_9 ;
wire \top/processor/sha_core/n12236_9 ;
wire \top/processor/sha_core/n12237_9 ;
wire \top/processor/sha_core/n12238_9 ;
wire \top/processor/sha_core/n12239_9 ;
wire \top/processor/sha_core/n12240_9 ;
wire \top/processor/sha_core/n12241_9 ;
wire \top/processor/sha_core/n12242_9 ;
wire \top/processor/sha_core/n12243_9 ;
wire \top/processor/sha_core/n12244_9 ;
wire \top/processor/sha_core/n12245_9 ;
wire \top/processor/sha_core/n12246_9 ;
wire \top/processor/sha_core/n12247_9 ;
wire \top/processor/sha_core/n12248_9 ;
wire \top/processor/sha_core/n12249_9 ;
wire \top/processor/sha_core/n12250_9 ;
wire \top/processor/sha_core/n12251_9 ;
wire \top/processor/sha_core/n12252_9 ;
wire \top/processor/sha_core/n12253_9 ;
wire \top/processor/sha_core/n12254_9 ;
wire \top/processor/sha_core/n12255_9 ;
wire \top/processor/sha_core/n12256_9 ;
wire \top/processor/sha_core/n12257_9 ;
wire \top/processor/sha_core/n12258_9 ;
wire \top/processor/sha_core/n12259_9 ;
wire \top/processor/sha_core/n12260_9 ;
wire \top/processor/sha_core/n12261_9 ;
wire \top/processor/sha_core/n12262_9 ;
wire \top/processor/sha_core/n12263_9 ;
wire \top/processor/sha_core/n12264_9 ;
wire \top/processor/sha_core/n12265_9 ;
wire \top/processor/sha_core/n12266_9 ;
wire \top/processor/sha_core/n12267_9 ;
wire \top/processor/sha_core/n12268_9 ;
wire \top/processor/sha_core/n12269_9 ;
wire \top/processor/sha_core/n12270_9 ;
wire \top/processor/sha_core/n12271_9 ;
wire \top/processor/sha_core/n12272_9 ;
wire \top/processor/sha_core/n12273_9 ;
wire \top/processor/sha_core/n12274_9 ;
wire \top/processor/sha_core/n12275_9 ;
wire \top/processor/sha_core/n12276_9 ;
wire \top/processor/sha_core/n12277_9 ;
wire \top/processor/sha_core/n12278_9 ;
wire \top/processor/sha_core/n12279_9 ;
wire \top/processor/sha_core/n12280_9 ;
wire \top/processor/sha_core/n12281_9 ;
wire \top/processor/sha_core/n12282_9 ;
wire \top/processor/sha_core/n12283_9 ;
wire \top/processor/sha_core/n12284_9 ;
wire \top/processor/sha_core/n12285_9 ;
wire \top/processor/sha_core/n12286_9 ;
wire \top/processor/sha_core/n12287_9 ;
wire \top/processor/sha_core/n12288_9 ;
wire \top/processor/sha_core/n12289_9 ;
wire \top/processor/sha_core/n12290_9 ;
wire \top/processor/sha_core/n12291_9 ;
wire \top/processor/sha_core/n12292_9 ;
wire \top/processor/sha_core/n12293_9 ;
wire \top/processor/sha_core/n12294_9 ;
wire \top/processor/sha_core/n12295_9 ;
wire \top/processor/sha_core/n12296_9 ;
wire \top/processor/sha_core/n12297_9 ;
wire \top/processor/sha_core/n12298_9 ;
wire \top/processor/sha_core/n12299_9 ;
wire \top/processor/sha_core/n12300_9 ;
wire \top/processor/sha_core/n12301_9 ;
wire \top/processor/sha_core/n12302_9 ;
wire \top/processor/sha_core/n12303_9 ;
wire \top/processor/sha_core/n12304_9 ;
wire \top/processor/sha_core/n12305_9 ;
wire \top/processor/sha_core/n12306_9 ;
wire \top/processor/sha_core/n12307_9 ;
wire \top/processor/sha_core/n12308_9 ;
wire \top/processor/sha_core/n12309_9 ;
wire \top/processor/sha_core/n12310_9 ;
wire \top/processor/sha_core/n12311_9 ;
wire \top/processor/sha_core/n12312_9 ;
wire \top/processor/sha_core/n12313_9 ;
wire \top/processor/sha_core/n12314_9 ;
wire \top/processor/sha_core/n12315_9 ;
wire \top/processor/sha_core/n12316_9 ;
wire \top/processor/sha_core/n12317_9 ;
wire \top/processor/sha_core/n12318_9 ;
wire \top/processor/sha_core/n12319_9 ;
wire \top/processor/sha_core/n12320_9 ;
wire \top/processor/sha_core/n12321_9 ;
wire \top/processor/sha_core/n12322_9 ;
wire \top/processor/sha_core/n12323_9 ;
wire \top/processor/sha_core/n12324_9 ;
wire \top/processor/sha_core/n12325_9 ;
wire \top/processor/sha_core/n12326_9 ;
wire \top/processor/sha_core/n12327_9 ;
wire \top/processor/sha_core/n12328_9 ;
wire \top/processor/sha_core/n12329_9 ;
wire \top/processor/sha_core/n12330_9 ;
wire \top/processor/sha_core/n12331_9 ;
wire \top/processor/sha_core/n12332_9 ;
wire \top/processor/sha_core/n12333_9 ;
wire \top/processor/sha_core/n12334_9 ;
wire \top/processor/sha_core/n12335_9 ;
wire \top/processor/sha_core/n12336_9 ;
wire \top/processor/sha_core/n12337_9 ;
wire \top/processor/sha_core/n12338_9 ;
wire \top/processor/sha_core/n12339_9 ;
wire \top/processor/sha_core/n12340_9 ;
wire \top/processor/sha_core/n12341_9 ;
wire \top/processor/sha_core/n12342_9 ;
wire \top/processor/sha_core/n12343_9 ;
wire \top/processor/sha_core/n12344_9 ;
wire \top/processor/sha_core/n12345_9 ;
wire \top/processor/sha_core/n12346_9 ;
wire \top/processor/sha_core/n12347_9 ;
wire \top/processor/sha_core/n12348_9 ;
wire \top/processor/sha_core/n12349_9 ;
wire \top/processor/sha_core/n12350_9 ;
wire \top/processor/sha_core/n12351_9 ;
wire \top/processor/sha_core/n12352_9 ;
wire \top/processor/sha_core/n12353_9 ;
wire \top/processor/sha_core/n12354_9 ;
wire \top/processor/sha_core/n12355_9 ;
wire \top/processor/sha_core/n12356_9 ;
wire \top/processor/sha_core/n12357_9 ;
wire \top/processor/sha_core/n12358_9 ;
wire \top/processor/sha_core/n12359_9 ;
wire \top/processor/sha_core/n12360_9 ;
wire \top/processor/sha_core/n12361_9 ;
wire \top/processor/sha_core/n12362_9 ;
wire \top/processor/sha_core/n12363_9 ;
wire \top/processor/sha_core/n12364_9 ;
wire \top/processor/sha_core/n12365_9 ;
wire \top/processor/sha_core/n12366_9 ;
wire \top/processor/sha_core/n12367_9 ;
wire \top/processor/sha_core/n12368_9 ;
wire \top/processor/sha_core/n12369_9 ;
wire \top/processor/sha_core/n12370_9 ;
wire \top/processor/sha_core/n12371_9 ;
wire \top/processor/sha_core/n12372_9 ;
wire \top/processor/sha_core/n12373_9 ;
wire \top/processor/sha_core/n12374_9 ;
wire \top/processor/sha_core/n12375_9 ;
wire \top/processor/sha_core/n12376_9 ;
wire \top/processor/sha_core/n12377_9 ;
wire \top/processor/sha_core/n12378_9 ;
wire \top/processor/sha_core/n12379_9 ;
wire \top/processor/sha_core/n12380_9 ;
wire \top/processor/sha_core/n12381_9 ;
wire \top/processor/sha_core/n12382_9 ;
wire \top/processor/sha_core/n12383_9 ;
wire \top/processor/sha_core/n12384_9 ;
wire \top/processor/sha_core/n12385_9 ;
wire \top/processor/sha_core/n12386_9 ;
wire \top/processor/sha_core/n12387_9 ;
wire \top/processor/sha_core/n12388_9 ;
wire \top/processor/sha_core/n12389_9 ;
wire \top/processor/sha_core/n12390_9 ;
wire \top/processor/sha_core/n11613_8 ;
wire \top/processor/sha_core/t_6_8 ;
wire \top/processor/sha_core/msg_idx_6_7 ;
wire \top/processor/sha_core/h0_31_8 ;
wire \top/processor/sha_core/w[2]_31_8 ;
wire \top/processor/sha_core/w[3]_31_8 ;
wire \top/processor/sha_core/w[4]_31_8 ;
wire \top/processor/sha_core/w[5]_31_8 ;
wire \top/processor/sha_core/w[6]_31_8 ;
wire \top/processor/sha_core/w[7]_31_8 ;
wire \top/processor/sha_core/w[8]_31_8 ;
wire \top/processor/sha_core/w[9]_31_8 ;
wire \top/processor/sha_core/w[10]_31_8 ;
wire \top/processor/sha_core/w[11]_31_8 ;
wire \top/processor/sha_core/w[12]_31_8 ;
wire \top/processor/sha_core/w[13]_31_8 ;
wire \top/processor/sha_core/w[14]_31_8 ;
wire \top/processor/sha_core/w[15]_31_8 ;
wire \top/processor/sha_core/w[16]_31_8 ;
wire \top/processor/sha_core/w[17]_31_8 ;
wire \top/processor/sha_core/w[18]_31_8 ;
wire \top/processor/sha_core/w[19]_31_8 ;
wire \top/processor/sha_core/w[20]_31_8 ;
wire \top/processor/sha_core/w[21]_31_8 ;
wire \top/processor/sha_core/w[22]_31_8 ;
wire \top/processor/sha_core/w[23]_31_8 ;
wire \top/processor/sha_core/w[24]_31_8 ;
wire \top/processor/sha_core/w[25]_31_8 ;
wire \top/processor/sha_core/w[26]_31_8 ;
wire \top/processor/sha_core/w[27]_31_8 ;
wire \top/processor/sha_core/w[28]_31_8 ;
wire \top/processor/sha_core/w[29]_31_8 ;
wire \top/processor/sha_core/w[30]_31_8 ;
wire \top/processor/sha_core/w[31]_31_8 ;
wire \top/processor/sha_core/w[48]_31_8 ;
wire \top/processor/sha_core/w[49]_31_8 ;
wire \top/processor/sha_core/w[50]_31_8 ;
wire \top/processor/sha_core/w[51]_31_8 ;
wire \top/processor/sha_core/w[52]_31_8 ;
wire \top/processor/sha_core/w[53]_31_8 ;
wire \top/processor/sha_core/w[54]_31_8 ;
wire \top/processor/sha_core/w[55]_31_8 ;
wire \top/processor/sha_core/w[56]_31_8 ;
wire \top/processor/sha_core/w[57]_31_8 ;
wire \top/processor/sha_core/w[58]_31_8 ;
wire \top/processor/sha_core/w[59]_31_8 ;
wire \top/processor/sha_core/w[60]_31_8 ;
wire \top/processor/sha_core/w[61]_31_8 ;
wire \top/processor/sha_core/w[62]_31_8 ;
wire \top/processor/sha_core/w[63]_31_8 ;
wire \top/processor/sha_core/h_31_8 ;
wire \top/processor/sha_core/n3453_7 ;
wire \top/processor/sha_core/n3452_7 ;
wire \top/processor/sha_core/n327_225 ;
wire \top/processor/sha_core/n328_225 ;
wire \top/processor/sha_core/n329_225 ;
wire \top/processor/sha_core/n330_225 ;
wire \top/processor/sha_core/n331_225 ;
wire \top/processor/sha_core/n332_225 ;
wire \top/processor/sha_core/n333_225 ;
wire \top/processor/sha_core/n334_225 ;
wire \top/processor/sha_core/n335_225 ;
wire \top/processor/sha_core/n336_225 ;
wire \top/processor/sha_core/n337_225 ;
wire \top/processor/sha_core/n338_225 ;
wire \top/processor/sha_core/n339_225 ;
wire \top/processor/sha_core/n340_225 ;
wire \top/processor/sha_core/n341_225 ;
wire \top/processor/sha_core/n342_225 ;
wire \top/processor/sha_core/n343_225 ;
wire \top/processor/sha_core/n344_225 ;
wire \top/processor/sha_core/n345_225 ;
wire \top/processor/sha_core/n346_225 ;
wire \top/processor/sha_core/n347_225 ;
wire \top/processor/sha_core/n348_225 ;
wire \top/processor/sha_core/n349_225 ;
wire \top/processor/sha_core/n350_225 ;
wire \top/processor/sha_core/n351_225 ;
wire \top/processor/sha_core/n352_225 ;
wire \top/processor/sha_core/n353_225 ;
wire \top/processor/sha_core/n354_225 ;
wire \top/processor/sha_core/n355_225 ;
wire \top/processor/sha_core/n356_225 ;
wire \top/processor/sha_core/n357_225 ;
wire \top/processor/sha_core/n358_225 ;
wire \top/processor/sha_core/n3607_187 ;
wire \top/processor/sha_core/n3607_189 ;
wire \top/processor/sha_core/n3607_191 ;
wire \top/processor/sha_core/n3607_193 ;
wire \top/processor/sha_core/n3608_187 ;
wire \top/processor/sha_core/n3608_189 ;
wire \top/processor/sha_core/n3608_191 ;
wire \top/processor/sha_core/n3608_193 ;
wire \top/processor/sha_core/n3609_187 ;
wire \top/processor/sha_core/n3609_189 ;
wire \top/processor/sha_core/n3609_191 ;
wire \top/processor/sha_core/n3609_193 ;
wire \top/processor/sha_core/n3610_187 ;
wire \top/processor/sha_core/n3610_189 ;
wire \top/processor/sha_core/n3610_191 ;
wire \top/processor/sha_core/n3610_193 ;
wire \top/processor/sha_core/n3611_187 ;
wire \top/processor/sha_core/n3611_189 ;
wire \top/processor/sha_core/n3611_191 ;
wire \top/processor/sha_core/n3611_193 ;
wire \top/processor/sha_core/n3612_187 ;
wire \top/processor/sha_core/n3612_189 ;
wire \top/processor/sha_core/n3612_191 ;
wire \top/processor/sha_core/n3612_193 ;
wire \top/processor/sha_core/n3613_187 ;
wire \top/processor/sha_core/n3613_189 ;
wire \top/processor/sha_core/n3613_191 ;
wire \top/processor/sha_core/n3613_193 ;
wire \top/processor/sha_core/n3614_187 ;
wire \top/processor/sha_core/n3614_189 ;
wire \top/processor/sha_core/n3614_191 ;
wire \top/processor/sha_core/n3614_193 ;
wire \top/processor/sha_core/n3615_187 ;
wire \top/processor/sha_core/n3615_189 ;
wire \top/processor/sha_core/n3615_191 ;
wire \top/processor/sha_core/n3615_193 ;
wire \top/processor/sha_core/n3616_187 ;
wire \top/processor/sha_core/n3616_189 ;
wire \top/processor/sha_core/n3616_191 ;
wire \top/processor/sha_core/n3616_193 ;
wire \top/processor/sha_core/n3617_187 ;
wire \top/processor/sha_core/n3617_189 ;
wire \top/processor/sha_core/n3617_191 ;
wire \top/processor/sha_core/n3617_193 ;
wire \top/processor/sha_core/n3618_187 ;
wire \top/processor/sha_core/n3618_189 ;
wire \top/processor/sha_core/n3618_191 ;
wire \top/processor/sha_core/n3618_193 ;
wire \top/processor/sha_core/n3619_187 ;
wire \top/processor/sha_core/n3619_189 ;
wire \top/processor/sha_core/n3619_191 ;
wire \top/processor/sha_core/n3619_193 ;
wire \top/processor/sha_core/n3620_187 ;
wire \top/processor/sha_core/n3620_189 ;
wire \top/processor/sha_core/n3620_191 ;
wire \top/processor/sha_core/n3620_193 ;
wire \top/processor/sha_core/n3621_187 ;
wire \top/processor/sha_core/n3621_189 ;
wire \top/processor/sha_core/n3621_191 ;
wire \top/processor/sha_core/n3621_193 ;
wire \top/processor/sha_core/n3622_187 ;
wire \top/processor/sha_core/n3622_189 ;
wire \top/processor/sha_core/n3622_191 ;
wire \top/processor/sha_core/n3622_193 ;
wire \top/processor/sha_core/n3623_187 ;
wire \top/processor/sha_core/n3623_189 ;
wire \top/processor/sha_core/n3623_191 ;
wire \top/processor/sha_core/n3623_193 ;
wire \top/processor/sha_core/n3624_187 ;
wire \top/processor/sha_core/n3624_189 ;
wire \top/processor/sha_core/n3624_191 ;
wire \top/processor/sha_core/n3624_193 ;
wire \top/processor/sha_core/n3625_187 ;
wire \top/processor/sha_core/n3625_189 ;
wire \top/processor/sha_core/n3625_191 ;
wire \top/processor/sha_core/n3625_193 ;
wire \top/processor/sha_core/n3626_187 ;
wire \top/processor/sha_core/n3626_189 ;
wire \top/processor/sha_core/n3626_191 ;
wire \top/processor/sha_core/n3626_193 ;
wire \top/processor/sha_core/n3627_187 ;
wire \top/processor/sha_core/n3627_189 ;
wire \top/processor/sha_core/n3627_191 ;
wire \top/processor/sha_core/n3627_193 ;
wire \top/processor/sha_core/n3628_187 ;
wire \top/processor/sha_core/n3628_189 ;
wire \top/processor/sha_core/n3628_191 ;
wire \top/processor/sha_core/n3628_193 ;
wire \top/processor/sha_core/n3629_187 ;
wire \top/processor/sha_core/n3629_189 ;
wire \top/processor/sha_core/n3629_191 ;
wire \top/processor/sha_core/n3629_193 ;
wire \top/processor/sha_core/n3630_187 ;
wire \top/processor/sha_core/n3630_189 ;
wire \top/processor/sha_core/n3630_191 ;
wire \top/processor/sha_core/n3630_193 ;
wire \top/processor/sha_core/n3631_187 ;
wire \top/processor/sha_core/n3631_189 ;
wire \top/processor/sha_core/n3631_191 ;
wire \top/processor/sha_core/n3631_193 ;
wire \top/processor/sha_core/n3632_187 ;
wire \top/processor/sha_core/n3632_189 ;
wire \top/processor/sha_core/n3632_191 ;
wire \top/processor/sha_core/n3632_193 ;
wire \top/processor/sha_core/n3633_187 ;
wire \top/processor/sha_core/n3633_189 ;
wire \top/processor/sha_core/n3633_191 ;
wire \top/processor/sha_core/n3633_193 ;
wire \top/processor/sha_core/n3634_187 ;
wire \top/processor/sha_core/n3634_189 ;
wire \top/processor/sha_core/n3634_191 ;
wire \top/processor/sha_core/n3634_193 ;
wire \top/processor/sha_core/n3635_187 ;
wire \top/processor/sha_core/n3635_189 ;
wire \top/processor/sha_core/n3635_191 ;
wire \top/processor/sha_core/n3635_193 ;
wire \top/processor/sha_core/n3636_187 ;
wire \top/processor/sha_core/n3636_189 ;
wire \top/processor/sha_core/n3636_191 ;
wire \top/processor/sha_core/n3636_193 ;
wire \top/processor/sha_core/n3637_187 ;
wire \top/processor/sha_core/n3637_189 ;
wire \top/processor/sha_core/n3637_191 ;
wire \top/processor/sha_core/n3637_193 ;
wire \top/processor/sha_core/n3638_187 ;
wire \top/processor/sha_core/n3638_189 ;
wire \top/processor/sha_core/n3638_191 ;
wire \top/processor/sha_core/n3638_193 ;
wire \top/processor/sha_core/n293_7162 ;
wire \top/processor/sha_core/n293_7164 ;
wire \top/processor/sha_core/n293_7166 ;
wire \top/processor/sha_core/n293_7168 ;
wire \top/processor/sha_core/n293_7170 ;
wire \top/processor/sha_core/n293_7172 ;
wire \top/processor/sha_core/n293_7174 ;
wire \top/processor/sha_core/n293_7176 ;
wire \top/processor/sha_core/n293_7178 ;
wire \top/processor/sha_core/n293_7180 ;
wire \top/processor/sha_core/n293_7182 ;
wire \top/processor/sha_core/n293_7184 ;
wire \top/processor/sha_core/n293_7186 ;
wire \top/processor/sha_core/n293_7188 ;
wire \top/processor/sha_core/n293_7190 ;
wire \top/processor/sha_core/n293_7192 ;
wire \top/processor/sha_core/n293_7194 ;
wire \top/processor/sha_core/n293_7196 ;
wire \top/processor/sha_core/n293_7198 ;
wire \top/processor/sha_core/n293_7200 ;
wire \top/processor/sha_core/n293_7202 ;
wire \top/processor/sha_core/n293_7204 ;
wire \top/processor/sha_core/n293_7206 ;
wire \top/processor/sha_core/n293_7208 ;
wire \top/processor/sha_core/n293_7210 ;
wire \top/processor/sha_core/n293_7212 ;
wire \top/processor/sha_core/n293_7214 ;
wire \top/processor/sha_core/n293_7216 ;
wire \top/processor/sha_core/n293_7218 ;
wire \top/processor/sha_core/n293_7220 ;
wire \top/processor/sha_core/n293_7222 ;
wire \top/processor/sha_core/n293_7224 ;
wire \top/processor/sha_core/n14445_10 ;
wire \top/processor/sha_core/n14442_9 ;
wire \top/processor/sha_core/n14440_9 ;
wire \top/processor/sha_core/n14439_9 ;
wire \top/processor/sha_core/n12134_11 ;
wire \top/processor/sha_core/n12133_11 ;
wire \top/processor/sha_core/n12132_11 ;
wire \top/processor/sha_core/n12131_11 ;
wire \top/processor/sha_core/n12130_11 ;
wire \top/processor/sha_core/n12129_11 ;
wire \top/processor/sha_core/n12128_11 ;
wire \top/processor/sha_core/n3462_11 ;
wire \top/processor/sha_core/n3461_11 ;
wire \top/processor/sha_core/n3460_11 ;
wire \top/processor/sha_core/n3459_9 ;
wire \top/processor/sha_core/n3578_11 ;
wire \top/processor/sha_core/n3834_9 ;
wire \top/processor/sha_core/n3766_4 ;
wire \top/processor/sha_core/n3766_5 ;
wire \top/processor/sha_core/n3767_4 ;
wire \top/processor/sha_core/n3767_5 ;
wire \top/processor/sha_core/n3768_4 ;
wire \top/processor/sha_core/n3768_5 ;
wire \top/processor/sha_core/n3769_4 ;
wire \top/processor/sha_core/n3769_5 ;
wire \top/processor/sha_core/n3769_6 ;
wire \top/processor/sha_core/n3770_4 ;
wire \top/processor/sha_core/n3770_5 ;
wire \top/processor/sha_core/n3771_4 ;
wire \top/processor/sha_core/n3771_5 ;
wire \top/processor/sha_core/n3772_4 ;
wire \top/processor/sha_core/n3772_5 ;
wire \top/processor/sha_core/n3773_4 ;
wire \top/processor/sha_core/n3773_5 ;
wire \top/processor/sha_core/n3774_4 ;
wire \top/processor/sha_core/n3774_5 ;
wire \top/processor/sha_core/n3775_4 ;
wire \top/processor/sha_core/n3775_5 ;
wire \top/processor/sha_core/n3776_4 ;
wire \top/processor/sha_core/n3776_5 ;
wire \top/processor/sha_core/n3777_4 ;
wire \top/processor/sha_core/n3778_4 ;
wire \top/processor/sha_core/n3779_4 ;
wire \top/processor/sha_core/n3780_4 ;
wire \top/processor/sha_core/n3781_4 ;
wire \top/processor/sha_core/n3782_4 ;
wire \top/processor/sha_core/n3783_4 ;
wire \top/processor/sha_core/n3784_4 ;
wire \top/processor/sha_core/n3785_4 ;
wire \top/processor/sha_core/n8430_4 ;
wire \top/processor/sha_core/n8430_5 ;
wire \top/processor/sha_core/n8430_6 ;
wire \top/processor/sha_core/n8431_4 ;
wire \top/processor/sha_core/n8431_5 ;
wire \top/processor/sha_core/n8432_4 ;
wire \top/processor/sha_core/n8432_5 ;
wire \top/processor/sha_core/n8433_4 ;
wire \top/processor/sha_core/n8433_5 ;
wire \top/processor/sha_core/n8434_4 ;
wire \top/processor/sha_core/n8434_5 ;
wire \top/processor/sha_core/n8435_4 ;
wire \top/processor/sha_core/n8435_5 ;
wire \top/processor/sha_core/n8436_4 ;
wire \top/processor/sha_core/n8436_5 ;
wire \top/processor/sha_core/n8437_4 ;
wire \top/processor/sha_core/n8437_5 ;
wire \top/processor/sha_core/n8438_4 ;
wire \top/processor/sha_core/n8438_5 ;
wire \top/processor/sha_core/n8439_4 ;
wire \top/processor/sha_core/n8440_4 ;
wire \top/processor/sha_core/n8440_5 ;
wire \top/processor/sha_core/n8441_4 ;
wire \top/processor/sha_core/n8441_5 ;
wire \top/processor/sha_core/n8442_4 ;
wire \top/processor/sha_core/n8443_4 ;
wire \top/processor/sha_core/n8443_5 ;
wire \top/processor/sha_core/n8444_4 ;
wire \top/processor/sha_core/n8444_5 ;
wire \top/processor/sha_core/n8445_4 ;
wire \top/processor/sha_core/n8445_5 ;
wire \top/processor/sha_core/n8446_4 ;
wire \top/processor/sha_core/n8446_5 ;
wire \top/processor/sha_core/n8447_4 ;
wire \top/processor/sha_core/n8447_5 ;
wire \top/processor/sha_core/n8448_4 ;
wire \top/processor/sha_core/n8448_5 ;
wire \top/processor/sha_core/n8449_4 ;
wire \top/processor/sha_core/n8449_5 ;
wire \top/processor/sha_core/n8450_4 ;
wire \top/processor/sha_core/n8451_4 ;
wire \top/processor/sha_core/n8451_5 ;
wire \top/processor/sha_core/n8452_4 ;
wire \top/processor/sha_core/n8452_5 ;
wire \top/processor/sha_core/n8453_4 ;
wire \top/processor/sha_core/n8453_5 ;
wire \top/processor/sha_core/n8454_4 ;
wire \top/processor/sha_core/n8454_5 ;
wire \top/processor/sha_core/n8455_4 ;
wire \top/processor/sha_core/n8455_5 ;
wire \top/processor/sha_core/n8456_4 ;
wire \top/processor/sha_core/n8456_5 ;
wire \top/processor/sha_core/n8457_4 ;
wire \top/processor/sha_core/n8458_4 ;
wire \top/processor/sha_core/n8458_5 ;
wire \top/processor/sha_core/n8459_4 ;
wire \top/processor/sha_core/n8459_5 ;
wire \top/processor/sha_core/n8460_4 ;
wire \top/processor/sha_core/n8460_5 ;
wire \top/processor/sha_core/n8461_4 ;
wire \top/processor/sha_core/n8461_5 ;
wire \top/processor/sha_core/state_0_9 ;
wire \top/processor/sha_core/w[0]_31_9 ;
wire \top/processor/sha_core/w[0]_31_10 ;
wire \top/processor/sha_core/w[1]_31_9 ;
wire \top/processor/sha_core/w[2]_31_9 ;
wire \top/processor/sha_core/w[3]_31_9 ;
wire \top/processor/sha_core/w[4]_31_9 ;
wire \top/processor/sha_core/w[5]_31_9 ;
wire \top/processor/sha_core/w[6]_31_9 ;
wire \top/processor/sha_core/w[8]_31_9 ;
wire \top/processor/sha_core/w[9]_31_9 ;
wire \top/processor/sha_core/w[10]_31_9 ;
wire \top/processor/sha_core/w[11]_31_9 ;
wire \top/processor/sha_core/w[12]_31_9 ;
wire \top/processor/sha_core/w[13]_31_9 ;
wire \top/processor/sha_core/w[14]_31_9 ;
wire \top/processor/sha_core/w[18]_31_9 ;
wire \top/processor/sha_core/w[19]_31_9 ;
wire \top/processor/sha_core/w[20]_31_9 ;
wire \top/processor/sha_core/w[21]_31_9 ;
wire \top/processor/sha_core/w[22]_31_9 ;
wire \top/processor/sha_core/w[40]_31_9 ;
wire \top/processor/sha_core/w[63]_31_9 ;
wire \top/processor/sha_core/n293_7225 ;
wire \top/processor/sha_core/n293_7226 ;
wire \top/processor/sha_core/n293_7227 ;
wire \top/processor/sha_core/n293_7228 ;
wire \top/processor/sha_core/n293_7229 ;
wire \top/processor/sha_core/n293_7230 ;
wire \top/processor/sha_core/n293_7231 ;
wire \top/processor/sha_core/n293_7232 ;
wire \top/processor/sha_core/n293_7233 ;
wire \top/processor/sha_core/n293_7235 ;
wire \top/processor/sha_core/n293_7236 ;
wire \top/processor/sha_core/n293_7237 ;
wire \top/processor/sha_core/n293_7238 ;
wire \top/processor/sha_core/n293_7239 ;
wire \top/processor/sha_core/n293_7240 ;
wire \top/processor/sha_core/n293_7241 ;
wire \top/processor/sha_core/n293_7242 ;
wire \top/processor/sha_core/n293_7243 ;
wire \top/processor/sha_core/n293_7244 ;
wire \top/processor/sha_core/n293_7245 ;
wire \top/processor/sha_core/n293_7246 ;
wire \top/processor/sha_core/n293_7247 ;
wire \top/processor/sha_core/n293_7248 ;
wire \top/processor/sha_core/n293_7249 ;
wire \top/processor/sha_core/n293_7250 ;
wire \top/processor/sha_core/n293_7251 ;
wire \top/processor/sha_core/n293_7252 ;
wire \top/processor/sha_core/n293_7253 ;
wire \top/processor/sha_core/n293_7254 ;
wire \top/processor/sha_core/n293_7255 ;
wire \top/processor/sha_core/n293_7256 ;
wire \top/processor/sha_core/n293_7257 ;
wire \top/processor/sha_core/n293_7258 ;
wire \top/processor/sha_core/n293_7259 ;
wire \top/processor/sha_core/n293_7260 ;
wire \top/processor/sha_core/n293_7261 ;
wire \top/processor/sha_core/n293_7262 ;
wire \top/processor/sha_core/n293_7263 ;
wire \top/processor/sha_core/n293_7264 ;
wire \top/processor/sha_core/n293_7265 ;
wire \top/processor/sha_core/n293_7266 ;
wire \top/processor/sha_core/n293_7267 ;
wire \top/processor/sha_core/n293_7268 ;
wire \top/processor/sha_core/n293_7269 ;
wire \top/processor/sha_core/n293_7270 ;
wire \top/processor/sha_core/n293_7271 ;
wire \top/processor/sha_core/n293_7272 ;
wire \top/processor/sha_core/n293_7273 ;
wire \top/processor/sha_core/n293_7274 ;
wire \top/processor/sha_core/n293_7275 ;
wire \top/processor/sha_core/n293_7276 ;
wire \top/processor/sha_core/n293_7277 ;
wire \top/processor/sha_core/n293_7278 ;
wire \top/processor/sha_core/n293_7279 ;
wire \top/processor/sha_core/n293_7280 ;
wire \top/processor/sha_core/n293_7281 ;
wire \top/processor/sha_core/n293_7282 ;
wire \top/processor/sha_core/n293_7283 ;
wire \top/processor/sha_core/n293_7284 ;
wire \top/processor/sha_core/n293_7285 ;
wire \top/processor/sha_core/n293_7286 ;
wire \top/processor/sha_core/n293_7287 ;
wire \top/processor/sha_core/n293_7288 ;
wire \top/processor/sha_core/n293_7289 ;
wire \top/processor/sha_core/n293_7290 ;
wire \top/processor/sha_core/n293_7291 ;
wire \top/processor/sha_core/n293_7292 ;
wire \top/processor/sha_core/n293_7293 ;
wire \top/processor/sha_core/n293_7294 ;
wire \top/processor/sha_core/n293_7295 ;
wire \top/processor/sha_core/n293_7296 ;
wire \top/processor/sha_core/n293_7297 ;
wire \top/processor/sha_core/n293_7298 ;
wire \top/processor/sha_core/n293_7299 ;
wire \top/processor/sha_core/n293_7300 ;
wire \top/processor/sha_core/n293_7301 ;
wire \top/processor/sha_core/n293_7302 ;
wire \top/processor/sha_core/n293_7303 ;
wire \top/processor/sha_core/n293_7304 ;
wire \top/processor/sha_core/n293_7305 ;
wire \top/processor/sha_core/n293_7306 ;
wire \top/processor/sha_core/n293_7307 ;
wire \top/processor/sha_core/n293_7308 ;
wire \top/processor/sha_core/n14441_10 ;
wire \top/processor/sha_core/n14439_10 ;
wire \top/processor/sha_core/n12131_12 ;
wire \top/processor/sha_core/n12129_12 ;
wire \top/processor/sha_core/n12128_12 ;
wire \top/processor/sha_core/n3578_12 ;
wire \top/processor/sha_core/n3766_6 ;
wire \top/processor/sha_core/n3766_7 ;
wire \top/processor/sha_core/n3766_8 ;
wire \top/processor/sha_core/n3766_9 ;
wire \top/processor/sha_core/n3766_10 ;
wire \top/processor/sha_core/n3767_6 ;
wire \top/processor/sha_core/n3767_7 ;
wire \top/processor/sha_core/n3767_8 ;
wire \top/processor/sha_core/n3767_9 ;
wire \top/processor/sha_core/n3768_6 ;
wire \top/processor/sha_core/n3768_7 ;
wire \top/processor/sha_core/n3768_8 ;
wire \top/processor/sha_core/n3768_9 ;
wire \top/processor/sha_core/n3769_7 ;
wire \top/processor/sha_core/n3769_8 ;
wire \top/processor/sha_core/n3769_9 ;
wire \top/processor/sha_core/n3769_10 ;
wire \top/processor/sha_core/n3769_11 ;
wire \top/processor/sha_core/n3769_12 ;
wire \top/processor/sha_core/n3770_6 ;
wire \top/processor/sha_core/n3770_7 ;
wire \top/processor/sha_core/n3770_8 ;
wire \top/processor/sha_core/n3770_9 ;
wire \top/processor/sha_core/n3771_6 ;
wire \top/processor/sha_core/n3771_7 ;
wire \top/processor/sha_core/n3771_8 ;
wire \top/processor/sha_core/n3771_9 ;
wire \top/processor/sha_core/n3772_6 ;
wire \top/processor/sha_core/n3772_7 ;
wire \top/processor/sha_core/n3772_8 ;
wire \top/processor/sha_core/n3772_9 ;
wire \top/processor/sha_core/n3773_6 ;
wire \top/processor/sha_core/n3773_7 ;
wire \top/processor/sha_core/n3773_8 ;
wire \top/processor/sha_core/n3773_9 ;
wire \top/processor/sha_core/n3774_6 ;
wire \top/processor/sha_core/n3774_7 ;
wire \top/processor/sha_core/n3774_8 ;
wire \top/processor/sha_core/n3774_9 ;
wire \top/processor/sha_core/n3775_6 ;
wire \top/processor/sha_core/n3775_7 ;
wire \top/processor/sha_core/n3775_8 ;
wire \top/processor/sha_core/n3775_9 ;
wire \top/processor/sha_core/n3776_6 ;
wire \top/processor/sha_core/n3776_7 ;
wire \top/processor/sha_core/n3776_8 ;
wire \top/processor/sha_core/n3776_9 ;
wire \top/processor/sha_core/n3777_5 ;
wire \top/processor/sha_core/n3777_6 ;
wire \top/processor/sha_core/n3778_5 ;
wire \top/processor/sha_core/n3778_6 ;
wire \top/processor/sha_core/n3779_5 ;
wire \top/processor/sha_core/n3779_6 ;
wire \top/processor/sha_core/n3780_5 ;
wire \top/processor/sha_core/n3780_6 ;
wire \top/processor/sha_core/n3781_5 ;
wire \top/processor/sha_core/n3781_6 ;
wire \top/processor/sha_core/n3782_5 ;
wire \top/processor/sha_core/n3782_6 ;
wire \top/processor/sha_core/n3783_5 ;
wire \top/processor/sha_core/n3783_6 ;
wire \top/processor/sha_core/n3784_5 ;
wire \top/processor/sha_core/n3784_6 ;
wire \top/processor/sha_core/n3785_5 ;
wire \top/processor/sha_core/n3785_6 ;
wire \top/processor/sha_core/n8430_7 ;
wire \top/processor/sha_core/n8430_8 ;
wire \top/processor/sha_core/n8430_9 ;
wire \top/processor/sha_core/n8430_10 ;
wire \top/processor/sha_core/n8430_11 ;
wire \top/processor/sha_core/n8430_12 ;
wire \top/processor/sha_core/n8430_13 ;
wire \top/processor/sha_core/n8431_6 ;
wire \top/processor/sha_core/n8431_7 ;
wire \top/processor/sha_core/n8431_8 ;
wire \top/processor/sha_core/n8431_9 ;
wire \top/processor/sha_core/n8431_10 ;
wire \top/processor/sha_core/n8431_11 ;
wire \top/processor/sha_core/n8431_12 ;
wire \top/processor/sha_core/n8432_6 ;
wire \top/processor/sha_core/n8432_7 ;
wire \top/processor/sha_core/n8432_8 ;
wire \top/processor/sha_core/n8432_9 ;
wire \top/processor/sha_core/n8432_10 ;
wire \top/processor/sha_core/n8432_11 ;
wire \top/processor/sha_core/n8433_6 ;
wire \top/processor/sha_core/n8433_7 ;
wire \top/processor/sha_core/n8433_8 ;
wire \top/processor/sha_core/n8433_9 ;
wire \top/processor/sha_core/n8433_10 ;
wire \top/processor/sha_core/n8433_11 ;
wire \top/processor/sha_core/n8434_6 ;
wire \top/processor/sha_core/n8434_7 ;
wire \top/processor/sha_core/n8434_8 ;
wire \top/processor/sha_core/n8434_9 ;
wire \top/processor/sha_core/n8434_10 ;
wire \top/processor/sha_core/n8434_11 ;
wire \top/processor/sha_core/n8435_6 ;
wire \top/processor/sha_core/n8435_7 ;
wire \top/processor/sha_core/n8435_8 ;
wire \top/processor/sha_core/n8435_9 ;
wire \top/processor/sha_core/n8435_10 ;
wire \top/processor/sha_core/n8435_11 ;
wire \top/processor/sha_core/n8435_12 ;
wire \top/processor/sha_core/n8435_13 ;
wire \top/processor/sha_core/n8436_6 ;
wire \top/processor/sha_core/n8436_7 ;
wire \top/processor/sha_core/n8436_8 ;
wire \top/processor/sha_core/n8436_9 ;
wire \top/processor/sha_core/n8436_10 ;
wire \top/processor/sha_core/n8436_11 ;
wire \top/processor/sha_core/n8437_6 ;
wire \top/processor/sha_core/n8437_7 ;
wire \top/processor/sha_core/n8437_8 ;
wire \top/processor/sha_core/n8437_9 ;
wire \top/processor/sha_core/n8437_10 ;
wire \top/processor/sha_core/n8437_11 ;
wire \top/processor/sha_core/n8438_6 ;
wire \top/processor/sha_core/n8438_7 ;
wire \top/processor/sha_core/n8438_8 ;
wire \top/processor/sha_core/n8438_9 ;
wire \top/processor/sha_core/n8438_10 ;
wire \top/processor/sha_core/n8438_11 ;
wire \top/processor/sha_core/n8439_5 ;
wire \top/processor/sha_core/n8439_6 ;
wire \top/processor/sha_core/n8440_6 ;
wire \top/processor/sha_core/n8440_7 ;
wire \top/processor/sha_core/n8440_8 ;
wire \top/processor/sha_core/n8440_9 ;
wire \top/processor/sha_core/n8440_10 ;
wire \top/processor/sha_core/n8440_11 ;
wire \top/processor/sha_core/n8441_6 ;
wire \top/processor/sha_core/n8441_7 ;
wire \top/processor/sha_core/n8441_8 ;
wire \top/processor/sha_core/n8441_9 ;
wire \top/processor/sha_core/n8441_10 ;
wire \top/processor/sha_core/n8441_11 ;
wire \top/processor/sha_core/n8442_5 ;
wire \top/processor/sha_core/n8442_6 ;
wire \top/processor/sha_core/n8442_7 ;
wire \top/processor/sha_core/n8442_8 ;
wire \top/processor/sha_core/n8443_6 ;
wire \top/processor/sha_core/n8443_7 ;
wire \top/processor/sha_core/n8443_8 ;
wire \top/processor/sha_core/n8443_9 ;
wire \top/processor/sha_core/n8443_10 ;
wire \top/processor/sha_core/n8443_11 ;
wire \top/processor/sha_core/n8444_6 ;
wire \top/processor/sha_core/n8444_7 ;
wire \top/processor/sha_core/n8444_8 ;
wire \top/processor/sha_core/n8444_9 ;
wire \top/processor/sha_core/n8444_10 ;
wire \top/processor/sha_core/n8444_11 ;
wire \top/processor/sha_core/n8445_6 ;
wire \top/processor/sha_core/n8445_7 ;
wire \top/processor/sha_core/n8445_8 ;
wire \top/processor/sha_core/n8445_9 ;
wire \top/processor/sha_core/n8445_10 ;
wire \top/processor/sha_core/n8445_11 ;
wire \top/processor/sha_core/n8445_12 ;
wire \top/processor/sha_core/n8445_13 ;
wire \top/processor/sha_core/n8446_6 ;
wire \top/processor/sha_core/n8446_7 ;
wire \top/processor/sha_core/n8446_8 ;
wire \top/processor/sha_core/n8446_9 ;
wire \top/processor/sha_core/n8446_10 ;
wire \top/processor/sha_core/n8446_11 ;
wire \top/processor/sha_core/n8447_6 ;
wire \top/processor/sha_core/n8447_7 ;
wire \top/processor/sha_core/n8447_8 ;
wire \top/processor/sha_core/n8447_9 ;
wire \top/processor/sha_core/n8447_10 ;
wire \top/processor/sha_core/n8447_11 ;
wire \top/processor/sha_core/n8448_6 ;
wire \top/processor/sha_core/n8448_7 ;
wire \top/processor/sha_core/n8448_8 ;
wire \top/processor/sha_core/n8448_9 ;
wire \top/processor/sha_core/n8448_10 ;
wire \top/processor/sha_core/n8448_11 ;
wire \top/processor/sha_core/n8449_6 ;
wire \top/processor/sha_core/n8449_7 ;
wire \top/processor/sha_core/n8449_8 ;
wire \top/processor/sha_core/n8449_9 ;
wire \top/processor/sha_core/n8449_10 ;
wire \top/processor/sha_core/n8449_11 ;
wire \top/processor/sha_core/n8450_5 ;
wire \top/processor/sha_core/n8450_6 ;
wire \top/processor/sha_core/n8450_7 ;
wire \top/processor/sha_core/n8450_8 ;
wire \top/processor/sha_core/n8451_6 ;
wire \top/processor/sha_core/n8451_7 ;
wire \top/processor/sha_core/n8451_8 ;
wire \top/processor/sha_core/n8451_9 ;
wire \top/processor/sha_core/n8451_10 ;
wire \top/processor/sha_core/n8451_11 ;
wire \top/processor/sha_core/n8451_12 ;
wire \top/processor/sha_core/n8451_13 ;
wire \top/processor/sha_core/n8452_6 ;
wire \top/processor/sha_core/n8452_7 ;
wire \top/processor/sha_core/n8452_8 ;
wire \top/processor/sha_core/n8452_9 ;
wire \top/processor/sha_core/n8452_10 ;
wire \top/processor/sha_core/n8452_11 ;
wire \top/processor/sha_core/n8453_6 ;
wire \top/processor/sha_core/n8453_7 ;
wire \top/processor/sha_core/n8453_8 ;
wire \top/processor/sha_core/n8453_9 ;
wire \top/processor/sha_core/n8453_10 ;
wire \top/processor/sha_core/n8453_11 ;
wire \top/processor/sha_core/n8454_6 ;
wire \top/processor/sha_core/n8454_7 ;
wire \top/processor/sha_core/n8454_8 ;
wire \top/processor/sha_core/n8454_9 ;
wire \top/processor/sha_core/n8454_10 ;
wire \top/processor/sha_core/n8454_11 ;
wire \top/processor/sha_core/n8455_6 ;
wire \top/processor/sha_core/n8455_7 ;
wire \top/processor/sha_core/n8455_8 ;
wire \top/processor/sha_core/n8455_9 ;
wire \top/processor/sha_core/n8455_10 ;
wire \top/processor/sha_core/n8455_11 ;
wire \top/processor/sha_core/n8455_12 ;
wire \top/processor/sha_core/n8455_13 ;
wire \top/processor/sha_core/n8456_6 ;
wire \top/processor/sha_core/n8456_7 ;
wire \top/processor/sha_core/n8456_8 ;
wire \top/processor/sha_core/n8456_9 ;
wire \top/processor/sha_core/n8456_10 ;
wire \top/processor/sha_core/n8456_11 ;
wire \top/processor/sha_core/n8457_5 ;
wire \top/processor/sha_core/n8457_6 ;
wire \top/processor/sha_core/n8458_6 ;
wire \top/processor/sha_core/n8458_7 ;
wire \top/processor/sha_core/n8458_8 ;
wire \top/processor/sha_core/n8458_9 ;
wire \top/processor/sha_core/n8458_10 ;
wire \top/processor/sha_core/n8458_11 ;
wire \top/processor/sha_core/n8459_6 ;
wire \top/processor/sha_core/n8459_7 ;
wire \top/processor/sha_core/n8459_8 ;
wire \top/processor/sha_core/n8459_9 ;
wire \top/processor/sha_core/n8459_10 ;
wire \top/processor/sha_core/n8459_11 ;
wire \top/processor/sha_core/n8460_6 ;
wire \top/processor/sha_core/n8460_7 ;
wire \top/processor/sha_core/n8460_8 ;
wire \top/processor/sha_core/n8460_9 ;
wire \top/processor/sha_core/n8460_10 ;
wire \top/processor/sha_core/n8460_11 ;
wire \top/processor/sha_core/n8461_6 ;
wire \top/processor/sha_core/n8461_7 ;
wire \top/processor/sha_core/n8461_8 ;
wire \top/processor/sha_core/n8461_9 ;
wire \top/processor/sha_core/n8461_10 ;
wire \top/processor/sha_core/n8461_11 ;
wire \top/processor/sha_core/n293_7309 ;
wire \top/processor/sha_core/n293_7310 ;
wire \top/processor/sha_core/n293_7311 ;
wire \top/processor/sha_core/n293_7312 ;
wire \top/processor/sha_core/n293_7313 ;
wire \top/processor/sha_core/n293_7314 ;
wire \top/processor/sha_core/n293_7315 ;
wire \top/processor/sha_core/n293_7316 ;
wire \top/processor/sha_core/n293_7317 ;
wire \top/processor/sha_core/n293_7318 ;
wire \top/processor/sha_core/n293_7319 ;
wire \top/processor/sha_core/n293_7320 ;
wire \top/processor/sha_core/n293_7322 ;
wire \top/processor/sha_core/n293_7324 ;
wire \top/processor/sha_core/n293_7325 ;
wire \top/processor/sha_core/n293_7326 ;
wire \top/processor/sha_core/n293_7327 ;
wire \top/processor/sha_core/n293_7328 ;
wire \top/processor/sha_core/n293_7329 ;
wire \top/processor/sha_core/n293_7330 ;
wire \top/processor/sha_core/n293_7331 ;
wire \top/processor/sha_core/n293_7332 ;
wire \top/processor/sha_core/n293_7333 ;
wire \top/processor/sha_core/n293_7334 ;
wire \top/processor/sha_core/n293_7335 ;
wire \top/processor/sha_core/n293_7336 ;
wire \top/processor/sha_core/n293_7337 ;
wire \top/processor/sha_core/n293_7338 ;
wire \top/processor/sha_core/n293_7339 ;
wire \top/processor/sha_core/n293_7340 ;
wire \top/processor/sha_core/n293_7341 ;
wire \top/processor/sha_core/n293_7342 ;
wire \top/processor/sha_core/n293_7343 ;
wire \top/processor/sha_core/n293_7344 ;
wire \top/processor/sha_core/n293_7345 ;
wire \top/processor/sha_core/n293_7346 ;
wire \top/processor/sha_core/n293_7347 ;
wire \top/processor/sha_core/n293_7348 ;
wire \top/processor/sha_core/n293_7349 ;
wire \top/processor/sha_core/n293_7350 ;
wire \top/processor/sha_core/n293_7351 ;
wire \top/processor/sha_core/n293_7352 ;
wire \top/processor/sha_core/n293_7353 ;
wire \top/processor/sha_core/n293_7354 ;
wire \top/processor/sha_core/n293_7355 ;
wire \top/processor/sha_core/n293_7356 ;
wire \top/processor/sha_core/n293_7357 ;
wire \top/processor/sha_core/n293_7358 ;
wire \top/processor/sha_core/n293_7359 ;
wire \top/processor/sha_core/n293_7360 ;
wire \top/processor/sha_core/n293_7361 ;
wire \top/processor/sha_core/n293_7362 ;
wire \top/processor/sha_core/n293_7363 ;
wire \top/processor/sha_core/n293_7364 ;
wire \top/processor/sha_core/n293_7365 ;
wire \top/processor/sha_core/n293_7366 ;
wire \top/processor/sha_core/n293_7367 ;
wire \top/processor/sha_core/n293_7368 ;
wire \top/processor/sha_core/n293_7369 ;
wire \top/processor/sha_core/n293_7370 ;
wire \top/processor/sha_core/n293_7371 ;
wire \top/processor/sha_core/n293_7372 ;
wire \top/processor/sha_core/n293_7373 ;
wire \top/processor/sha_core/n293_7374 ;
wire \top/processor/sha_core/n293_7375 ;
wire \top/processor/sha_core/n293_7376 ;
wire \top/processor/sha_core/n293_7377 ;
wire \top/processor/sha_core/n293_7378 ;
wire \top/processor/sha_core/n293_7379 ;
wire \top/processor/sha_core/n293_7380 ;
wire \top/processor/sha_core/n293_7381 ;
wire \top/processor/sha_core/n293_7382 ;
wire \top/processor/sha_core/n293_7383 ;
wire \top/processor/sha_core/n3766_11 ;
wire \top/processor/sha_core/n3766_12 ;
wire \top/processor/sha_core/n3766_13 ;
wire \top/processor/sha_core/n3766_14 ;
wire \top/processor/sha_core/n3767_10 ;
wire \top/processor/sha_core/n3767_11 ;
wire \top/processor/sha_core/n3767_12 ;
wire \top/processor/sha_core/n3767_13 ;
wire \top/processor/sha_core/n3768_10 ;
wire \top/processor/sha_core/n3768_11 ;
wire \top/processor/sha_core/n3768_12 ;
wire \top/processor/sha_core/n3768_13 ;
wire \top/processor/sha_core/n3769_13 ;
wire \top/processor/sha_core/n3769_14 ;
wire \top/processor/sha_core/n3769_15 ;
wire \top/processor/sha_core/n3769_16 ;
wire \top/processor/sha_core/n3769_17 ;
wire \top/processor/sha_core/n3769_18 ;
wire \top/processor/sha_core/n3770_10 ;
wire \top/processor/sha_core/n3770_11 ;
wire \top/processor/sha_core/n3770_12 ;
wire \top/processor/sha_core/n3770_13 ;
wire \top/processor/sha_core/n3771_10 ;
wire \top/processor/sha_core/n3771_11 ;
wire \top/processor/sha_core/n3771_12 ;
wire \top/processor/sha_core/n3771_13 ;
wire \top/processor/sha_core/n3772_10 ;
wire \top/processor/sha_core/n3772_11 ;
wire \top/processor/sha_core/n3772_12 ;
wire \top/processor/sha_core/n3772_13 ;
wire \top/processor/sha_core/n3773_10 ;
wire \top/processor/sha_core/n3773_11 ;
wire \top/processor/sha_core/n3773_12 ;
wire \top/processor/sha_core/n3773_13 ;
wire \top/processor/sha_core/n3774_10 ;
wire \top/processor/sha_core/n3774_11 ;
wire \top/processor/sha_core/n3774_12 ;
wire \top/processor/sha_core/n3774_13 ;
wire \top/processor/sha_core/n3775_10 ;
wire \top/processor/sha_core/n3775_11 ;
wire \top/processor/sha_core/n3775_12 ;
wire \top/processor/sha_core/n3775_13 ;
wire \top/processor/sha_core/n3776_10 ;
wire \top/processor/sha_core/n3776_11 ;
wire \top/processor/sha_core/n3776_12 ;
wire \top/processor/sha_core/n3776_13 ;
wire \top/processor/sha_core/n3777_7 ;
wire \top/processor/sha_core/n3777_8 ;
wire \top/processor/sha_core/n3778_7 ;
wire \top/processor/sha_core/n3778_8 ;
wire \top/processor/sha_core/n3779_7 ;
wire \top/processor/sha_core/n3779_8 ;
wire \top/processor/sha_core/n3780_7 ;
wire \top/processor/sha_core/n3780_8 ;
wire \top/processor/sha_core/n3781_7 ;
wire \top/processor/sha_core/n3781_8 ;
wire \top/processor/sha_core/n3782_7 ;
wire \top/processor/sha_core/n3782_8 ;
wire \top/processor/sha_core/n3783_7 ;
wire \top/processor/sha_core/n3783_8 ;
wire \top/processor/sha_core/n3784_7 ;
wire \top/processor/sha_core/n3784_8 ;
wire \top/processor/sha_core/n3785_7 ;
wire \top/processor/sha_core/n3785_8 ;
wire \top/processor/sha_core/n8430_14 ;
wire \top/processor/sha_core/n8430_15 ;
wire \top/processor/sha_core/n8431_13 ;
wire \top/processor/sha_core/n8431_14 ;
wire \top/processor/sha_core/n8432_12 ;
wire \top/processor/sha_core/n8432_13 ;
wire \top/processor/sha_core/n8433_12 ;
wire \top/processor/sha_core/n8433_13 ;
wire \top/processor/sha_core/n8434_12 ;
wire \top/processor/sha_core/n8434_13 ;
wire \top/processor/sha_core/n8436_12 ;
wire \top/processor/sha_core/n8436_13 ;
wire \top/processor/sha_core/n8437_12 ;
wire \top/processor/sha_core/n8437_13 ;
wire \top/processor/sha_core/n8438_12 ;
wire \top/processor/sha_core/n8438_13 ;
wire \top/processor/sha_core/n8439_7 ;
wire \top/processor/sha_core/n8439_8 ;
wire \top/processor/sha_core/n8439_9 ;
wire \top/processor/sha_core/n8439_10 ;
wire \top/processor/sha_core/n8439_11 ;
wire \top/processor/sha_core/n8439_12 ;
wire \top/processor/sha_core/n8440_12 ;
wire \top/processor/sha_core/n8440_13 ;
wire \top/processor/sha_core/n8441_12 ;
wire \top/processor/sha_core/n8441_13 ;
wire \top/processor/sha_core/n8442_9 ;
wire \top/processor/sha_core/n8442_10 ;
wire \top/processor/sha_core/n8442_11 ;
wire \top/processor/sha_core/n8442_12 ;
wire \top/processor/sha_core/n8442_13 ;
wire \top/processor/sha_core/n8443_12 ;
wire \top/processor/sha_core/n8443_13 ;
wire \top/processor/sha_core/n8444_12 ;
wire \top/processor/sha_core/n8444_13 ;
wire \top/processor/sha_core/n8446_12 ;
wire \top/processor/sha_core/n8446_13 ;
wire \top/processor/sha_core/n8447_12 ;
wire \top/processor/sha_core/n8447_13 ;
wire \top/processor/sha_core/n8448_12 ;
wire \top/processor/sha_core/n8448_13 ;
wire \top/processor/sha_core/n8449_12 ;
wire \top/processor/sha_core/n8449_13 ;
wire \top/processor/sha_core/n8450_9 ;
wire \top/processor/sha_core/n8450_10 ;
wire \top/processor/sha_core/n8450_11 ;
wire \top/processor/sha_core/n8450_12 ;
wire \top/processor/sha_core/n8450_13 ;
wire \top/processor/sha_core/n8452_12 ;
wire \top/processor/sha_core/n8452_13 ;
wire \top/processor/sha_core/n8453_12 ;
wire \top/processor/sha_core/n8453_13 ;
wire \top/processor/sha_core/n8454_12 ;
wire \top/processor/sha_core/n8454_13 ;
wire \top/processor/sha_core/n8456_12 ;
wire \top/processor/sha_core/n8456_13 ;
wire \top/processor/sha_core/n8457_7 ;
wire \top/processor/sha_core/n8457_8 ;
wire \top/processor/sha_core/n8457_9 ;
wire \top/processor/sha_core/n8457_10 ;
wire \top/processor/sha_core/n8457_11 ;
wire \top/processor/sha_core/n8458_12 ;
wire \top/processor/sha_core/n8458_13 ;
wire \top/processor/sha_core/n8459_12 ;
wire \top/processor/sha_core/n8459_13 ;
wire \top/processor/sha_core/n8460_12 ;
wire \top/processor/sha_core/n8460_13 ;
wire \top/processor/sha_core/n8461_12 ;
wire \top/processor/sha_core/n8461_13 ;
wire \top/processor/sha_core/n8439_13 ;
wire \top/processor/sha_core/n8439_14 ;
wire \top/processor/sha_core/n8442_14 ;
wire \top/processor/sha_core/n8450_14 ;
wire \top/processor/sha_core/n8457_12 ;
wire \top/processor/sha_core/n8457_13 ;
wire \top/processor/sha_core/n8457_14 ;
wire \top/processor/sha_core/n293_7386 ;
wire \top/processor/sha_core/n293_7388 ;
wire \top/processor/sha_core/n3766_16 ;
wire \top/processor/sha_core/n3767_15 ;
wire \top/processor/sha_core/n3768_15 ;
wire \top/processor/sha_core/n3607_196 ;
wire \top/processor/sha_core/w[31]_31_11 ;
wire \top/processor/sha_core/w[23]_31_11 ;
wire \top/processor/sha_core/w[15]_31_11 ;
wire \top/processor/sha_core/w[7]_31_11 ;
wire \top/processor/sha_core/w[2]_31_12 ;
wire \top/processor/sha_core/w[47]_31_10 ;
wire \top/processor/sha_core/w[46]_31_10 ;
wire \top/processor/sha_core/w[45]_31_10 ;
wire \top/processor/sha_core/w[44]_31_10 ;
wire \top/processor/sha_core/w[43]_31_10 ;
wire \top/processor/sha_core/w[42]_31_10 ;
wire \top/processor/sha_core/w[41]_31_10 ;
wire \top/processor/sha_core/w[40]_31_11 ;
wire \top/processor/sha_core/n3577_11 ;
wire \top/processor/sha_core/w[39]_31_10 ;
wire \top/processor/sha_core/w[38]_31_10 ;
wire \top/processor/sha_core/w[37]_31_10 ;
wire \top/processor/sha_core/w[36]_31_10 ;
wire \top/processor/sha_core/w[35]_31_10 ;
wire \top/processor/sha_core/w[34]_31_10 ;
wire \top/processor/sha_core/w[33]_31_10 ;
wire \top/processor/sha_core/w[32]_31_10 ;
wire \top/processor/sha_core/w[1]_31_11 ;
wire \top/processor/sha_core/w[0]_31_12 ;
wire \top/processor/sha_core/n14441_12 ;
wire \top/processor/sha_core/n14443_11 ;
wire \top/processor/sha_core/n14444_11 ;
wire \top/processor/sha_core/n3544_5 ;
wire \top/processor/sha_core/n3542_5 ;
wire \top/processor/sha_core/n11871_15 ;
wire \top/processor/sha_core/n11870_15 ;
wire \top/processor/sha_core/n3924_1 ;
wire \top/processor/sha_core/n3924_2 ;
wire \top/processor/sha_core/n3923_1 ;
wire \top/processor/sha_core/n3923_2 ;
wire \top/processor/sha_core/n3922_1 ;
wire \top/processor/sha_core/n3922_2 ;
wire \top/processor/sha_core/n3921_1 ;
wire \top/processor/sha_core/n3921_2 ;
wire \top/processor/sha_core/n3920_1 ;
wire \top/processor/sha_core/n3920_2 ;
wire \top/processor/sha_core/n3919_1 ;
wire \top/processor/sha_core/n3919_2 ;
wire \top/processor/sha_core/n3918_1 ;
wire \top/processor/sha_core/n3918_2 ;
wire \top/processor/sha_core/n3917_1 ;
wire \top/processor/sha_core/n3917_2 ;
wire \top/processor/sha_core/n3916_1 ;
wire \top/processor/sha_core/n3916_2 ;
wire \top/processor/sha_core/n3915_1 ;
wire \top/processor/sha_core/n3915_2 ;
wire \top/processor/sha_core/n3914_1 ;
wire \top/processor/sha_core/n3914_2 ;
wire \top/processor/sha_core/n3913_1 ;
wire \top/processor/sha_core/n3913_2 ;
wire \top/processor/sha_core/n3912_1 ;
wire \top/processor/sha_core/n3912_2 ;
wire \top/processor/sha_core/n3911_1 ;
wire \top/processor/sha_core/n3911_2 ;
wire \top/processor/sha_core/n3910_1 ;
wire \top/processor/sha_core/n3910_2 ;
wire \top/processor/sha_core/n3909_1 ;
wire \top/processor/sha_core/n3909_2 ;
wire \top/processor/sha_core/n3908_1 ;
wire \top/processor/sha_core/n3908_2 ;
wire \top/processor/sha_core/n3907_1 ;
wire \top/processor/sha_core/n3907_2 ;
wire \top/processor/sha_core/n3906_1 ;
wire \top/processor/sha_core/n3906_2 ;
wire \top/processor/sha_core/n3905_1 ;
wire \top/processor/sha_core/n3905_2 ;
wire \top/processor/sha_core/n3904_1 ;
wire \top/processor/sha_core/n3904_2 ;
wire \top/processor/sha_core/n3903_1 ;
wire \top/processor/sha_core/n3903_2 ;
wire \top/processor/sha_core/n3902_1 ;
wire \top/processor/sha_core/n3902_2 ;
wire \top/processor/sha_core/n3901_1 ;
wire \top/processor/sha_core/n3901_2 ;
wire \top/processor/sha_core/n3900_1 ;
wire \top/processor/sha_core/n3900_2 ;
wire \top/processor/sha_core/n3899_1 ;
wire \top/processor/sha_core/n3899_2 ;
wire \top/processor/sha_core/n3898_1 ;
wire \top/processor/sha_core/n3898_2 ;
wire \top/processor/sha_core/n3897_1 ;
wire \top/processor/sha_core/n3897_2 ;
wire \top/processor/sha_core/n3896_1 ;
wire \top/processor/sha_core/n3896_2 ;
wire \top/processor/sha_core/n3895_1 ;
wire \top/processor/sha_core/n3895_2 ;
wire \top/processor/sha_core/n3894_1 ;
wire \top/processor/sha_core/n3894_2 ;
wire \top/processor/sha_core/n3893_1 ;
wire \top/processor/sha_core/n3893_0_COUT ;
wire \top/processor/sha_core/n3924_3 ;
wire \top/processor/sha_core/n3924_4 ;
wire \top/processor/sha_core/n3923_3 ;
wire \top/processor/sha_core/n3923_4 ;
wire \top/processor/sha_core/n3922_3 ;
wire \top/processor/sha_core/n3922_4 ;
wire \top/processor/sha_core/n3921_3 ;
wire \top/processor/sha_core/n3921_4 ;
wire \top/processor/sha_core/n3920_3 ;
wire \top/processor/sha_core/n3920_4 ;
wire \top/processor/sha_core/n3919_3 ;
wire \top/processor/sha_core/n3919_4 ;
wire \top/processor/sha_core/n3918_3 ;
wire \top/processor/sha_core/n3918_4 ;
wire \top/processor/sha_core/n3917_3 ;
wire \top/processor/sha_core/n3917_4 ;
wire \top/processor/sha_core/n3916_3 ;
wire \top/processor/sha_core/n3916_4 ;
wire \top/processor/sha_core/n3915_3 ;
wire \top/processor/sha_core/n3915_4 ;
wire \top/processor/sha_core/n3914_3 ;
wire \top/processor/sha_core/n3914_4 ;
wire \top/processor/sha_core/n3913_3 ;
wire \top/processor/sha_core/n3913_4 ;
wire \top/processor/sha_core/n3912_3 ;
wire \top/processor/sha_core/n3912_4 ;
wire \top/processor/sha_core/n3911_3 ;
wire \top/processor/sha_core/n3911_4 ;
wire \top/processor/sha_core/n3910_3 ;
wire \top/processor/sha_core/n3910_4 ;
wire \top/processor/sha_core/n3909_3 ;
wire \top/processor/sha_core/n3909_4 ;
wire \top/processor/sha_core/n3908_3 ;
wire \top/processor/sha_core/n3908_4 ;
wire \top/processor/sha_core/n3907_3 ;
wire \top/processor/sha_core/n3907_4 ;
wire \top/processor/sha_core/n3906_3 ;
wire \top/processor/sha_core/n3906_4 ;
wire \top/processor/sha_core/n3905_3 ;
wire \top/processor/sha_core/n3905_4 ;
wire \top/processor/sha_core/n3904_3 ;
wire \top/processor/sha_core/n3904_4 ;
wire \top/processor/sha_core/n3903_3 ;
wire \top/processor/sha_core/n3903_4 ;
wire \top/processor/sha_core/n3902_3 ;
wire \top/processor/sha_core/n3902_4 ;
wire \top/processor/sha_core/n3901_3 ;
wire \top/processor/sha_core/n3901_4 ;
wire \top/processor/sha_core/n3900_3 ;
wire \top/processor/sha_core/n3900_4 ;
wire \top/processor/sha_core/n3899_3 ;
wire \top/processor/sha_core/n3899_4 ;
wire \top/processor/sha_core/n3898_3 ;
wire \top/processor/sha_core/n3898_4 ;
wire \top/processor/sha_core/n3897_3 ;
wire \top/processor/sha_core/n3897_4 ;
wire \top/processor/sha_core/n3896_3 ;
wire \top/processor/sha_core/n3896_4 ;
wire \top/processor/sha_core/n3895_3 ;
wire \top/processor/sha_core/n3895_4 ;
wire \top/processor/sha_core/n3894_3 ;
wire \top/processor/sha_core/n3894_4 ;
wire \top/processor/sha_core/n3893_3 ;
wire \top/processor/sha_core/n3893_1_COUT ;
wire \top/processor/sha_core/n3924_5 ;
wire \top/processor/sha_core/n3924_6 ;
wire \top/processor/sha_core/n3923_5 ;
wire \top/processor/sha_core/n3923_6 ;
wire \top/processor/sha_core/n3922_5 ;
wire \top/processor/sha_core/n3922_6 ;
wire \top/processor/sha_core/n3921_5 ;
wire \top/processor/sha_core/n3921_6 ;
wire \top/processor/sha_core/n3920_5 ;
wire \top/processor/sha_core/n3920_6 ;
wire \top/processor/sha_core/n3919_5 ;
wire \top/processor/sha_core/n3919_6 ;
wire \top/processor/sha_core/n3918_5 ;
wire \top/processor/sha_core/n3918_6 ;
wire \top/processor/sha_core/n3917_5 ;
wire \top/processor/sha_core/n3917_6 ;
wire \top/processor/sha_core/n3916_5 ;
wire \top/processor/sha_core/n3916_6 ;
wire \top/processor/sha_core/n3915_5 ;
wire \top/processor/sha_core/n3915_6 ;
wire \top/processor/sha_core/n3914_5 ;
wire \top/processor/sha_core/n3914_6 ;
wire \top/processor/sha_core/n3913_5 ;
wire \top/processor/sha_core/n3913_6 ;
wire \top/processor/sha_core/n3912_5 ;
wire \top/processor/sha_core/n3912_6 ;
wire \top/processor/sha_core/n3911_5 ;
wire \top/processor/sha_core/n3911_6 ;
wire \top/processor/sha_core/n3910_5 ;
wire \top/processor/sha_core/n3910_6 ;
wire \top/processor/sha_core/n3909_5 ;
wire \top/processor/sha_core/n3909_6 ;
wire \top/processor/sha_core/n3908_5 ;
wire \top/processor/sha_core/n3908_6 ;
wire \top/processor/sha_core/n3907_5 ;
wire \top/processor/sha_core/n3907_6 ;
wire \top/processor/sha_core/n3906_5 ;
wire \top/processor/sha_core/n3906_6 ;
wire \top/processor/sha_core/n3905_5 ;
wire \top/processor/sha_core/n3905_6 ;
wire \top/processor/sha_core/n3904_5 ;
wire \top/processor/sha_core/n3904_6 ;
wire \top/processor/sha_core/n3903_5 ;
wire \top/processor/sha_core/n3903_6 ;
wire \top/processor/sha_core/n3902_5 ;
wire \top/processor/sha_core/n3902_6 ;
wire \top/processor/sha_core/n3901_5 ;
wire \top/processor/sha_core/n3901_6 ;
wire \top/processor/sha_core/n3900_5 ;
wire \top/processor/sha_core/n3900_6 ;
wire \top/processor/sha_core/n3899_5 ;
wire \top/processor/sha_core/n3899_6 ;
wire \top/processor/sha_core/n3898_5 ;
wire \top/processor/sha_core/n3898_6 ;
wire \top/processor/sha_core/n3897_5 ;
wire \top/processor/sha_core/n3897_6 ;
wire \top/processor/sha_core/n3896_5 ;
wire \top/processor/sha_core/n3896_6 ;
wire \top/processor/sha_core/n3895_5 ;
wire \top/processor/sha_core/n3895_6 ;
wire \top/processor/sha_core/n3894_5 ;
wire \top/processor/sha_core/n3894_6 ;
wire \top/processor/sha_core/n3893_5 ;
wire \top/processor/sha_core/n3893_2_COUT ;
wire \top/processor/sha_core/n10857_1 ;
wire \top/processor/sha_core/n10857_2 ;
wire \top/processor/sha_core/n10856_1 ;
wire \top/processor/sha_core/n10856_2 ;
wire \top/processor/sha_core/n10855_1 ;
wire \top/processor/sha_core/n10855_2 ;
wire \top/processor/sha_core/n10854_1 ;
wire \top/processor/sha_core/n10854_2 ;
wire \top/processor/sha_core/n10853_1 ;
wire \top/processor/sha_core/n10853_2 ;
wire \top/processor/sha_core/n10852_1 ;
wire \top/processor/sha_core/n10852_2 ;
wire \top/processor/sha_core/n10851_1 ;
wire \top/processor/sha_core/n10851_2 ;
wire \top/processor/sha_core/n10850_1 ;
wire \top/processor/sha_core/n10850_2 ;
wire \top/processor/sha_core/n10849_1 ;
wire \top/processor/sha_core/n10849_2 ;
wire \top/processor/sha_core/n10848_1 ;
wire \top/processor/sha_core/n10848_2 ;
wire \top/processor/sha_core/n10847_1 ;
wire \top/processor/sha_core/n10847_2 ;
wire \top/processor/sha_core/n10846_1 ;
wire \top/processor/sha_core/n10846_2 ;
wire \top/processor/sha_core/n10845_1 ;
wire \top/processor/sha_core/n10845_2 ;
wire \top/processor/sha_core/n10844_1 ;
wire \top/processor/sha_core/n10844_2 ;
wire \top/processor/sha_core/n10843_1 ;
wire \top/processor/sha_core/n10843_2 ;
wire \top/processor/sha_core/n10842_1 ;
wire \top/processor/sha_core/n10842_2 ;
wire \top/processor/sha_core/n10841_1 ;
wire \top/processor/sha_core/n10841_2 ;
wire \top/processor/sha_core/n10840_1 ;
wire \top/processor/sha_core/n10840_2 ;
wire \top/processor/sha_core/n10839_1 ;
wire \top/processor/sha_core/n10839_2 ;
wire \top/processor/sha_core/n10838_1 ;
wire \top/processor/sha_core/n10838_2 ;
wire \top/processor/sha_core/n10837_1 ;
wire \top/processor/sha_core/n10837_2 ;
wire \top/processor/sha_core/n10836_1 ;
wire \top/processor/sha_core/n10836_2 ;
wire \top/processor/sha_core/n10835_1 ;
wire \top/processor/sha_core/n10835_2 ;
wire \top/processor/sha_core/n10834_1 ;
wire \top/processor/sha_core/n10834_2 ;
wire \top/processor/sha_core/n10833_1 ;
wire \top/processor/sha_core/n10833_2 ;
wire \top/processor/sha_core/n10832_1 ;
wire \top/processor/sha_core/n10832_2 ;
wire \top/processor/sha_core/n10831_1 ;
wire \top/processor/sha_core/n10831_2 ;
wire \top/processor/sha_core/n10830_1 ;
wire \top/processor/sha_core/n10830_2 ;
wire \top/processor/sha_core/n10829_1 ;
wire \top/processor/sha_core/n10829_2 ;
wire \top/processor/sha_core/n10828_1 ;
wire \top/processor/sha_core/n10828_2 ;
wire \top/processor/sha_core/n10827_1 ;
wire \top/processor/sha_core/n10827_2 ;
wire \top/processor/sha_core/n10826_1 ;
wire \top/processor/sha_core/n10826_0_COUT ;
wire \top/processor/sha_core/n10890_1 ;
wire \top/processor/sha_core/n10890_2 ;
wire \top/processor/sha_core/n10889_1 ;
wire \top/processor/sha_core/n10889_2 ;
wire \top/processor/sha_core/n10888_1 ;
wire \top/processor/sha_core/n10888_2 ;
wire \top/processor/sha_core/n10887_1 ;
wire \top/processor/sha_core/n10887_2 ;
wire \top/processor/sha_core/n10886_1 ;
wire \top/processor/sha_core/n10886_2 ;
wire \top/processor/sha_core/n10885_1 ;
wire \top/processor/sha_core/n10885_2 ;
wire \top/processor/sha_core/n10884_1 ;
wire \top/processor/sha_core/n10884_2 ;
wire \top/processor/sha_core/n10883_1 ;
wire \top/processor/sha_core/n10883_2 ;
wire \top/processor/sha_core/n10882_1 ;
wire \top/processor/sha_core/n10882_2 ;
wire \top/processor/sha_core/n10881_1 ;
wire \top/processor/sha_core/n10881_2 ;
wire \top/processor/sha_core/n10880_1 ;
wire \top/processor/sha_core/n10880_2 ;
wire \top/processor/sha_core/n10879_1 ;
wire \top/processor/sha_core/n10879_2 ;
wire \top/processor/sha_core/n10878_1 ;
wire \top/processor/sha_core/n10878_2 ;
wire \top/processor/sha_core/n10877_1 ;
wire \top/processor/sha_core/n10877_2 ;
wire \top/processor/sha_core/n10876_1 ;
wire \top/processor/sha_core/n10876_2 ;
wire \top/processor/sha_core/n10875_1 ;
wire \top/processor/sha_core/n10875_2 ;
wire \top/processor/sha_core/n10874_1 ;
wire \top/processor/sha_core/n10874_2 ;
wire \top/processor/sha_core/n10873_1 ;
wire \top/processor/sha_core/n10873_2 ;
wire \top/processor/sha_core/n10872_1 ;
wire \top/processor/sha_core/n10872_2 ;
wire \top/processor/sha_core/n10871_1 ;
wire \top/processor/sha_core/n10871_2 ;
wire \top/processor/sha_core/n10870_1 ;
wire \top/processor/sha_core/n10870_2 ;
wire \top/processor/sha_core/n10869_1 ;
wire \top/processor/sha_core/n10869_2 ;
wire \top/processor/sha_core/n10868_1 ;
wire \top/processor/sha_core/n10868_2 ;
wire \top/processor/sha_core/n10867_1 ;
wire \top/processor/sha_core/n10867_2 ;
wire \top/processor/sha_core/n10866_1 ;
wire \top/processor/sha_core/n10866_2 ;
wire \top/processor/sha_core/n10865_1 ;
wire \top/processor/sha_core/n10865_2 ;
wire \top/processor/sha_core/n10864_1 ;
wire \top/processor/sha_core/n10864_2 ;
wire \top/processor/sha_core/n10863_1 ;
wire \top/processor/sha_core/n10863_2 ;
wire \top/processor/sha_core/n10862_1 ;
wire \top/processor/sha_core/n10862_2 ;
wire \top/processor/sha_core/n10861_1 ;
wire \top/processor/sha_core/n10861_2 ;
wire \top/processor/sha_core/n10860_1 ;
wire \top/processor/sha_core/n10860_2 ;
wire \top/processor/sha_core/n10859_1 ;
wire \top/processor/sha_core/n10859_0_COUT ;
wire \top/processor/sha_core/n10923_1 ;
wire \top/processor/sha_core/n10923_2 ;
wire \top/processor/sha_core/n10922_1 ;
wire \top/processor/sha_core/n10922_2 ;
wire \top/processor/sha_core/n10921_1 ;
wire \top/processor/sha_core/n10921_2 ;
wire \top/processor/sha_core/n10920_1 ;
wire \top/processor/sha_core/n10920_2 ;
wire \top/processor/sha_core/n10919_1 ;
wire \top/processor/sha_core/n10919_2 ;
wire \top/processor/sha_core/n10918_1 ;
wire \top/processor/sha_core/n10918_2 ;
wire \top/processor/sha_core/n10917_1 ;
wire \top/processor/sha_core/n10917_2 ;
wire \top/processor/sha_core/n10916_1 ;
wire \top/processor/sha_core/n10916_2 ;
wire \top/processor/sha_core/n10915_1 ;
wire \top/processor/sha_core/n10915_2 ;
wire \top/processor/sha_core/n10914_1 ;
wire \top/processor/sha_core/n10914_2 ;
wire \top/processor/sha_core/n10913_1 ;
wire \top/processor/sha_core/n10913_2 ;
wire \top/processor/sha_core/n10912_1 ;
wire \top/processor/sha_core/n10912_2 ;
wire \top/processor/sha_core/n10911_1 ;
wire \top/processor/sha_core/n10911_2 ;
wire \top/processor/sha_core/n10910_1 ;
wire \top/processor/sha_core/n10910_2 ;
wire \top/processor/sha_core/n10909_1 ;
wire \top/processor/sha_core/n10909_2 ;
wire \top/processor/sha_core/n10908_1 ;
wire \top/processor/sha_core/n10908_2 ;
wire \top/processor/sha_core/n10907_1 ;
wire \top/processor/sha_core/n10907_2 ;
wire \top/processor/sha_core/n10906_1 ;
wire \top/processor/sha_core/n10906_2 ;
wire \top/processor/sha_core/n10905_1 ;
wire \top/processor/sha_core/n10905_2 ;
wire \top/processor/sha_core/n10904_1 ;
wire \top/processor/sha_core/n10904_2 ;
wire \top/processor/sha_core/n10903_1 ;
wire \top/processor/sha_core/n10903_2 ;
wire \top/processor/sha_core/n10902_1 ;
wire \top/processor/sha_core/n10902_2 ;
wire \top/processor/sha_core/n10901_1 ;
wire \top/processor/sha_core/n10901_2 ;
wire \top/processor/sha_core/n10900_1 ;
wire \top/processor/sha_core/n10900_2 ;
wire \top/processor/sha_core/n10899_1 ;
wire \top/processor/sha_core/n10899_2 ;
wire \top/processor/sha_core/n10898_1 ;
wire \top/processor/sha_core/n10898_2 ;
wire \top/processor/sha_core/n10897_1 ;
wire \top/processor/sha_core/n10897_2 ;
wire \top/processor/sha_core/n10896_1 ;
wire \top/processor/sha_core/n10896_2 ;
wire \top/processor/sha_core/n10895_1 ;
wire \top/processor/sha_core/n10895_2 ;
wire \top/processor/sha_core/n10894_1 ;
wire \top/processor/sha_core/n10894_2 ;
wire \top/processor/sha_core/n10893_1 ;
wire \top/processor/sha_core/n10893_2 ;
wire \top/processor/sha_core/n10892_1 ;
wire \top/processor/sha_core/n10892_0_COUT ;
wire \top/processor/sha_core/n10956_1 ;
wire \top/processor/sha_core/n10956_2 ;
wire \top/processor/sha_core/n10955_1 ;
wire \top/processor/sha_core/n10955_2 ;
wire \top/processor/sha_core/n10954_1 ;
wire \top/processor/sha_core/n10954_2 ;
wire \top/processor/sha_core/n10953_1 ;
wire \top/processor/sha_core/n10953_2 ;
wire \top/processor/sha_core/n10952_1 ;
wire \top/processor/sha_core/n10952_2 ;
wire \top/processor/sha_core/n10951_1 ;
wire \top/processor/sha_core/n10951_2 ;
wire \top/processor/sha_core/n10950_1 ;
wire \top/processor/sha_core/n10950_2 ;
wire \top/processor/sha_core/n10949_1 ;
wire \top/processor/sha_core/n10949_2 ;
wire \top/processor/sha_core/n10948_1 ;
wire \top/processor/sha_core/n10948_2 ;
wire \top/processor/sha_core/n10947_1 ;
wire \top/processor/sha_core/n10947_2 ;
wire \top/processor/sha_core/n10946_1 ;
wire \top/processor/sha_core/n10946_2 ;
wire \top/processor/sha_core/n10945_1 ;
wire \top/processor/sha_core/n10945_2 ;
wire \top/processor/sha_core/n10944_1 ;
wire \top/processor/sha_core/n10944_2 ;
wire \top/processor/sha_core/n10943_1 ;
wire \top/processor/sha_core/n10943_2 ;
wire \top/processor/sha_core/n10942_1 ;
wire \top/processor/sha_core/n10942_2 ;
wire \top/processor/sha_core/n10941_1 ;
wire \top/processor/sha_core/n10941_2 ;
wire \top/processor/sha_core/n10940_1 ;
wire \top/processor/sha_core/n10940_2 ;
wire \top/processor/sha_core/n10939_1 ;
wire \top/processor/sha_core/n10939_2 ;
wire \top/processor/sha_core/n10938_1 ;
wire \top/processor/sha_core/n10938_2 ;
wire \top/processor/sha_core/n10937_1 ;
wire \top/processor/sha_core/n10937_2 ;
wire \top/processor/sha_core/n10936_1 ;
wire \top/processor/sha_core/n10936_2 ;
wire \top/processor/sha_core/n10935_1 ;
wire \top/processor/sha_core/n10935_2 ;
wire \top/processor/sha_core/n10934_1 ;
wire \top/processor/sha_core/n10934_2 ;
wire \top/processor/sha_core/n10933_1 ;
wire \top/processor/sha_core/n10933_2 ;
wire \top/processor/sha_core/n10932_1 ;
wire \top/processor/sha_core/n10932_2 ;
wire \top/processor/sha_core/n10931_1 ;
wire \top/processor/sha_core/n10931_2 ;
wire \top/processor/sha_core/n10930_1 ;
wire \top/processor/sha_core/n10930_2 ;
wire \top/processor/sha_core/n10929_1 ;
wire \top/processor/sha_core/n10929_2 ;
wire \top/processor/sha_core/n10928_1 ;
wire \top/processor/sha_core/n10928_2 ;
wire \top/processor/sha_core/n10927_1 ;
wire \top/processor/sha_core/n10927_2 ;
wire \top/processor/sha_core/n10926_1 ;
wire \top/processor/sha_core/n10926_2 ;
wire \top/processor/sha_core/n10925_1 ;
wire \top/processor/sha_core/n10925_0_COUT ;
wire \top/processor/sha_core/n10989_1 ;
wire \top/processor/sha_core/n10989_2 ;
wire \top/processor/sha_core/n10988_1 ;
wire \top/processor/sha_core/n10988_2 ;
wire \top/processor/sha_core/n10987_1 ;
wire \top/processor/sha_core/n10987_2 ;
wire \top/processor/sha_core/n10986_1 ;
wire \top/processor/sha_core/n10986_2 ;
wire \top/processor/sha_core/n10985_1 ;
wire \top/processor/sha_core/n10985_2 ;
wire \top/processor/sha_core/n10984_1 ;
wire \top/processor/sha_core/n10984_2 ;
wire \top/processor/sha_core/n10983_1 ;
wire \top/processor/sha_core/n10983_2 ;
wire \top/processor/sha_core/n10982_1 ;
wire \top/processor/sha_core/n10982_2 ;
wire \top/processor/sha_core/n10981_1 ;
wire \top/processor/sha_core/n10981_2 ;
wire \top/processor/sha_core/n10980_1 ;
wire \top/processor/sha_core/n10980_2 ;
wire \top/processor/sha_core/n10979_1 ;
wire \top/processor/sha_core/n10979_2 ;
wire \top/processor/sha_core/n10978_1 ;
wire \top/processor/sha_core/n10978_2 ;
wire \top/processor/sha_core/n10977_1 ;
wire \top/processor/sha_core/n10977_2 ;
wire \top/processor/sha_core/n10976_1 ;
wire \top/processor/sha_core/n10976_2 ;
wire \top/processor/sha_core/n10975_1 ;
wire \top/processor/sha_core/n10975_2 ;
wire \top/processor/sha_core/n10974_1 ;
wire \top/processor/sha_core/n10974_2 ;
wire \top/processor/sha_core/n10973_1 ;
wire \top/processor/sha_core/n10973_2 ;
wire \top/processor/sha_core/n10972_1 ;
wire \top/processor/sha_core/n10972_2 ;
wire \top/processor/sha_core/n10971_1 ;
wire \top/processor/sha_core/n10971_2 ;
wire \top/processor/sha_core/n10970_1 ;
wire \top/processor/sha_core/n10970_2 ;
wire \top/processor/sha_core/n10969_1 ;
wire \top/processor/sha_core/n10969_2 ;
wire \top/processor/sha_core/n10968_1 ;
wire \top/processor/sha_core/n10968_2 ;
wire \top/processor/sha_core/n10967_1 ;
wire \top/processor/sha_core/n10967_2 ;
wire \top/processor/sha_core/n10966_1 ;
wire \top/processor/sha_core/n10966_2 ;
wire \top/processor/sha_core/n10965_1 ;
wire \top/processor/sha_core/n10965_2 ;
wire \top/processor/sha_core/n10964_1 ;
wire \top/processor/sha_core/n10964_2 ;
wire \top/processor/sha_core/n10963_1 ;
wire \top/processor/sha_core/n10963_2 ;
wire \top/processor/sha_core/n10962_1 ;
wire \top/processor/sha_core/n10962_2 ;
wire \top/processor/sha_core/n10961_1 ;
wire \top/processor/sha_core/n10961_2 ;
wire \top/processor/sha_core/n10960_1 ;
wire \top/processor/sha_core/n10960_2 ;
wire \top/processor/sha_core/n10959_1 ;
wire \top/processor/sha_core/n10959_2 ;
wire \top/processor/sha_core/n10958_1 ;
wire \top/processor/sha_core/n10958_0_COUT ;
wire \top/processor/sha_core/n11022_1 ;
wire \top/processor/sha_core/n11022_2 ;
wire \top/processor/sha_core/n11021_1 ;
wire \top/processor/sha_core/n11021_2 ;
wire \top/processor/sha_core/n11020_1 ;
wire \top/processor/sha_core/n11020_2 ;
wire \top/processor/sha_core/n11019_1 ;
wire \top/processor/sha_core/n11019_2 ;
wire \top/processor/sha_core/n11018_1 ;
wire \top/processor/sha_core/n11018_2 ;
wire \top/processor/sha_core/n11017_1 ;
wire \top/processor/sha_core/n11017_2 ;
wire \top/processor/sha_core/n11016_1 ;
wire \top/processor/sha_core/n11016_2 ;
wire \top/processor/sha_core/n11015_1 ;
wire \top/processor/sha_core/n11015_2 ;
wire \top/processor/sha_core/n11014_1 ;
wire \top/processor/sha_core/n11014_2 ;
wire \top/processor/sha_core/n11013_1 ;
wire \top/processor/sha_core/n11013_2 ;
wire \top/processor/sha_core/n11012_1 ;
wire \top/processor/sha_core/n11012_2 ;
wire \top/processor/sha_core/n11011_1 ;
wire \top/processor/sha_core/n11011_2 ;
wire \top/processor/sha_core/n11010_1 ;
wire \top/processor/sha_core/n11010_2 ;
wire \top/processor/sha_core/n11009_1 ;
wire \top/processor/sha_core/n11009_2 ;
wire \top/processor/sha_core/n11008_1 ;
wire \top/processor/sha_core/n11008_2 ;
wire \top/processor/sha_core/n11007_1 ;
wire \top/processor/sha_core/n11007_2 ;
wire \top/processor/sha_core/n11006_1 ;
wire \top/processor/sha_core/n11006_2 ;
wire \top/processor/sha_core/n11005_1 ;
wire \top/processor/sha_core/n11005_2 ;
wire \top/processor/sha_core/n11004_1 ;
wire \top/processor/sha_core/n11004_2 ;
wire \top/processor/sha_core/n11003_1 ;
wire \top/processor/sha_core/n11003_2 ;
wire \top/processor/sha_core/n11002_1 ;
wire \top/processor/sha_core/n11002_2 ;
wire \top/processor/sha_core/n11001_1 ;
wire \top/processor/sha_core/n11001_2 ;
wire \top/processor/sha_core/n11000_1 ;
wire \top/processor/sha_core/n11000_2 ;
wire \top/processor/sha_core/n10999_1 ;
wire \top/processor/sha_core/n10999_2 ;
wire \top/processor/sha_core/n10998_1 ;
wire \top/processor/sha_core/n10998_2 ;
wire \top/processor/sha_core/n10997_1 ;
wire \top/processor/sha_core/n10997_2 ;
wire \top/processor/sha_core/n10996_1 ;
wire \top/processor/sha_core/n10996_2 ;
wire \top/processor/sha_core/n10995_1 ;
wire \top/processor/sha_core/n10995_2 ;
wire \top/processor/sha_core/n10994_1 ;
wire \top/processor/sha_core/n10994_2 ;
wire \top/processor/sha_core/n10993_1 ;
wire \top/processor/sha_core/n10993_2 ;
wire \top/processor/sha_core/n10992_1 ;
wire \top/processor/sha_core/n10992_2 ;
wire \top/processor/sha_core/n10991_1 ;
wire \top/processor/sha_core/n10991_0_COUT ;
wire \top/processor/sha_core/n11055_1 ;
wire \top/processor/sha_core/n11055_2 ;
wire \top/processor/sha_core/n11054_1 ;
wire \top/processor/sha_core/n11054_2 ;
wire \top/processor/sha_core/n11053_1 ;
wire \top/processor/sha_core/n11053_2 ;
wire \top/processor/sha_core/n11052_1 ;
wire \top/processor/sha_core/n11052_2 ;
wire \top/processor/sha_core/n11051_1 ;
wire \top/processor/sha_core/n11051_2 ;
wire \top/processor/sha_core/n11050_1 ;
wire \top/processor/sha_core/n11050_2 ;
wire \top/processor/sha_core/n11049_1 ;
wire \top/processor/sha_core/n11049_2 ;
wire \top/processor/sha_core/n11048_1 ;
wire \top/processor/sha_core/n11048_2 ;
wire \top/processor/sha_core/n11047_1 ;
wire \top/processor/sha_core/n11047_2 ;
wire \top/processor/sha_core/n11046_1 ;
wire \top/processor/sha_core/n11046_2 ;
wire \top/processor/sha_core/n11045_1 ;
wire \top/processor/sha_core/n11045_2 ;
wire \top/processor/sha_core/n11044_1 ;
wire \top/processor/sha_core/n11044_2 ;
wire \top/processor/sha_core/n11043_1 ;
wire \top/processor/sha_core/n11043_2 ;
wire \top/processor/sha_core/n11042_1 ;
wire \top/processor/sha_core/n11042_2 ;
wire \top/processor/sha_core/n11041_1 ;
wire \top/processor/sha_core/n11041_2 ;
wire \top/processor/sha_core/n11040_1 ;
wire \top/processor/sha_core/n11040_2 ;
wire \top/processor/sha_core/n11039_1 ;
wire \top/processor/sha_core/n11039_2 ;
wire \top/processor/sha_core/n11038_1 ;
wire \top/processor/sha_core/n11038_2 ;
wire \top/processor/sha_core/n11037_1 ;
wire \top/processor/sha_core/n11037_2 ;
wire \top/processor/sha_core/n11036_1 ;
wire \top/processor/sha_core/n11036_2 ;
wire \top/processor/sha_core/n11035_1 ;
wire \top/processor/sha_core/n11035_2 ;
wire \top/processor/sha_core/n11034_1 ;
wire \top/processor/sha_core/n11034_2 ;
wire \top/processor/sha_core/n11033_1 ;
wire \top/processor/sha_core/n11033_2 ;
wire \top/processor/sha_core/n11032_1 ;
wire \top/processor/sha_core/n11032_2 ;
wire \top/processor/sha_core/n11031_1 ;
wire \top/processor/sha_core/n11031_2 ;
wire \top/processor/sha_core/n11030_1 ;
wire \top/processor/sha_core/n11030_2 ;
wire \top/processor/sha_core/n11029_1 ;
wire \top/processor/sha_core/n11029_2 ;
wire \top/processor/sha_core/n11028_1 ;
wire \top/processor/sha_core/n11028_2 ;
wire \top/processor/sha_core/n11027_1 ;
wire \top/processor/sha_core/n11027_2 ;
wire \top/processor/sha_core/n11026_1 ;
wire \top/processor/sha_core/n11026_2 ;
wire \top/processor/sha_core/n11025_1 ;
wire \top/processor/sha_core/n11025_2 ;
wire \top/processor/sha_core/n11024_1 ;
wire \top/processor/sha_core/n11024_0_COUT ;
wire \top/processor/sha_core/n11088_1 ;
wire \top/processor/sha_core/n11088_2 ;
wire \top/processor/sha_core/n11087_1 ;
wire \top/processor/sha_core/n11087_2 ;
wire \top/processor/sha_core/n11086_1 ;
wire \top/processor/sha_core/n11086_2 ;
wire \top/processor/sha_core/n11085_1 ;
wire \top/processor/sha_core/n11085_2 ;
wire \top/processor/sha_core/n11084_1 ;
wire \top/processor/sha_core/n11084_2 ;
wire \top/processor/sha_core/n11083_1 ;
wire \top/processor/sha_core/n11083_2 ;
wire \top/processor/sha_core/n11082_1 ;
wire \top/processor/sha_core/n11082_2 ;
wire \top/processor/sha_core/n11081_1 ;
wire \top/processor/sha_core/n11081_2 ;
wire \top/processor/sha_core/n11080_1 ;
wire \top/processor/sha_core/n11080_2 ;
wire \top/processor/sha_core/n11079_1 ;
wire \top/processor/sha_core/n11079_2 ;
wire \top/processor/sha_core/n11078_1 ;
wire \top/processor/sha_core/n11078_2 ;
wire \top/processor/sha_core/n11077_1 ;
wire \top/processor/sha_core/n11077_2 ;
wire \top/processor/sha_core/n11076_1 ;
wire \top/processor/sha_core/n11076_2 ;
wire \top/processor/sha_core/n11075_1 ;
wire \top/processor/sha_core/n11075_2 ;
wire \top/processor/sha_core/n11074_1 ;
wire \top/processor/sha_core/n11074_2 ;
wire \top/processor/sha_core/n11073_1 ;
wire \top/processor/sha_core/n11073_2 ;
wire \top/processor/sha_core/n11072_1 ;
wire \top/processor/sha_core/n11072_2 ;
wire \top/processor/sha_core/n11071_1 ;
wire \top/processor/sha_core/n11071_2 ;
wire \top/processor/sha_core/n11070_1 ;
wire \top/processor/sha_core/n11070_2 ;
wire \top/processor/sha_core/n11069_1 ;
wire \top/processor/sha_core/n11069_2 ;
wire \top/processor/sha_core/n11068_1 ;
wire \top/processor/sha_core/n11068_2 ;
wire \top/processor/sha_core/n11067_1 ;
wire \top/processor/sha_core/n11067_2 ;
wire \top/processor/sha_core/n11066_1 ;
wire \top/processor/sha_core/n11066_2 ;
wire \top/processor/sha_core/n11065_1 ;
wire \top/processor/sha_core/n11065_2 ;
wire \top/processor/sha_core/n11064_1 ;
wire \top/processor/sha_core/n11064_2 ;
wire \top/processor/sha_core/n11063_1 ;
wire \top/processor/sha_core/n11063_2 ;
wire \top/processor/sha_core/n11062_1 ;
wire \top/processor/sha_core/n11062_2 ;
wire \top/processor/sha_core/n11061_1 ;
wire \top/processor/sha_core/n11061_2 ;
wire \top/processor/sha_core/n11060_1 ;
wire \top/processor/sha_core/n11060_2 ;
wire \top/processor/sha_core/n11059_1 ;
wire \top/processor/sha_core/n11059_2 ;
wire \top/processor/sha_core/n11058_1 ;
wire \top/processor/sha_core/n11058_2 ;
wire \top/processor/sha_core/n11057_1 ;
wire \top/processor/sha_core/n11057_0_COUT ;
wire \top/processor/sha_core/n10783_3 ;
wire \top/processor/sha_core/n10783_4 ;
wire \top/processor/sha_core/n10782_3 ;
wire \top/processor/sha_core/n10782_4 ;
wire \top/processor/sha_core/n10781_3 ;
wire \top/processor/sha_core/n10781_4 ;
wire \top/processor/sha_core/n10780_3 ;
wire \top/processor/sha_core/n10780_4 ;
wire \top/processor/sha_core/n10779_3 ;
wire \top/processor/sha_core/n10779_4 ;
wire \top/processor/sha_core/n10778_3 ;
wire \top/processor/sha_core/n10778_4 ;
wire \top/processor/sha_core/n10777_3 ;
wire \top/processor/sha_core/n10777_4 ;
wire \top/processor/sha_core/n10776_3 ;
wire \top/processor/sha_core/n10776_4 ;
wire \top/processor/sha_core/n10775_3 ;
wire \top/processor/sha_core/n10775_4 ;
wire \top/processor/sha_core/n10774_3 ;
wire \top/processor/sha_core/n10774_4 ;
wire \top/processor/sha_core/n10773_3 ;
wire \top/processor/sha_core/n10773_4 ;
wire \top/processor/sha_core/n10772_3 ;
wire \top/processor/sha_core/n10772_4 ;
wire \top/processor/sha_core/n10771_3 ;
wire \top/processor/sha_core/n10771_4 ;
wire \top/processor/sha_core/n10770_3 ;
wire \top/processor/sha_core/n10770_4 ;
wire \top/processor/sha_core/n10769_3 ;
wire \top/processor/sha_core/n10769_4 ;
wire \top/processor/sha_core/n10768_3 ;
wire \top/processor/sha_core/n10768_4 ;
wire \top/processor/sha_core/n10767_3 ;
wire \top/processor/sha_core/n10767_4 ;
wire \top/processor/sha_core/n10766_3 ;
wire \top/processor/sha_core/n10766_4 ;
wire \top/processor/sha_core/n10765_3 ;
wire \top/processor/sha_core/n10765_4 ;
wire \top/processor/sha_core/n10764_3 ;
wire \top/processor/sha_core/n10764_4 ;
wire \top/processor/sha_core/n10763_3 ;
wire \top/processor/sha_core/n10763_4 ;
wire \top/processor/sha_core/n10762_3 ;
wire \top/processor/sha_core/n10762_4 ;
wire \top/processor/sha_core/n10761_3 ;
wire \top/processor/sha_core/n10761_4 ;
wire \top/processor/sha_core/n10760_3 ;
wire \top/processor/sha_core/n10760_4 ;
wire \top/processor/sha_core/n10759_3 ;
wire \top/processor/sha_core/n10759_4 ;
wire \top/processor/sha_core/n10758_3 ;
wire \top/processor/sha_core/n10758_4 ;
wire \top/processor/sha_core/n10757_3 ;
wire \top/processor/sha_core/n10757_4 ;
wire \top/processor/sha_core/n10756_3 ;
wire \top/processor/sha_core/n10756_4 ;
wire \top/processor/sha_core/n10755_3 ;
wire \top/processor/sha_core/n10755_4 ;
wire \top/processor/sha_core/n10754_3 ;
wire \top/processor/sha_core/n10754_4 ;
wire \top/processor/sha_core/n10753_3 ;
wire \top/processor/sha_core/n10753_4 ;
wire \top/processor/sha_core/n10752_3 ;
wire \top/processor/sha_core/n10752_0_COUT ;
wire \top/processor/sha_core/n10783_5 ;
wire \top/processor/sha_core/n10783_6 ;
wire \top/processor/sha_core/n10782_5 ;
wire \top/processor/sha_core/n10782_6 ;
wire \top/processor/sha_core/n10781_5 ;
wire \top/processor/sha_core/n10781_6 ;
wire \top/processor/sha_core/n10780_5 ;
wire \top/processor/sha_core/n10780_6 ;
wire \top/processor/sha_core/n10779_5 ;
wire \top/processor/sha_core/n10779_6 ;
wire \top/processor/sha_core/n10778_5 ;
wire \top/processor/sha_core/n10778_6 ;
wire \top/processor/sha_core/n10777_5 ;
wire \top/processor/sha_core/n10777_6 ;
wire \top/processor/sha_core/n10776_5 ;
wire \top/processor/sha_core/n10776_6 ;
wire \top/processor/sha_core/n10775_5 ;
wire \top/processor/sha_core/n10775_6 ;
wire \top/processor/sha_core/n10774_5 ;
wire \top/processor/sha_core/n10774_6 ;
wire \top/processor/sha_core/n10773_5 ;
wire \top/processor/sha_core/n10773_6 ;
wire \top/processor/sha_core/n10772_5 ;
wire \top/processor/sha_core/n10772_6 ;
wire \top/processor/sha_core/n10771_5 ;
wire \top/processor/sha_core/n10771_6 ;
wire \top/processor/sha_core/n10770_5 ;
wire \top/processor/sha_core/n10770_6 ;
wire \top/processor/sha_core/n10769_5 ;
wire \top/processor/sha_core/n10769_6 ;
wire \top/processor/sha_core/n10768_5 ;
wire \top/processor/sha_core/n10768_6 ;
wire \top/processor/sha_core/n10767_5 ;
wire \top/processor/sha_core/n10767_6 ;
wire \top/processor/sha_core/n10766_5 ;
wire \top/processor/sha_core/n10766_6 ;
wire \top/processor/sha_core/n10765_5 ;
wire \top/processor/sha_core/n10765_6 ;
wire \top/processor/sha_core/n10764_5 ;
wire \top/processor/sha_core/n10764_6 ;
wire \top/processor/sha_core/n10763_5 ;
wire \top/processor/sha_core/n10763_6 ;
wire \top/processor/sha_core/n10762_5 ;
wire \top/processor/sha_core/n10762_6 ;
wire \top/processor/sha_core/n10761_5 ;
wire \top/processor/sha_core/n10761_6 ;
wire \top/processor/sha_core/n10760_5 ;
wire \top/processor/sha_core/n10760_6 ;
wire \top/processor/sha_core/n10759_5 ;
wire \top/processor/sha_core/n10759_6 ;
wire \top/processor/sha_core/n10758_5 ;
wire \top/processor/sha_core/n10758_6 ;
wire \top/processor/sha_core/n10757_5 ;
wire \top/processor/sha_core/n10757_6 ;
wire \top/processor/sha_core/n10756_5 ;
wire \top/processor/sha_core/n10756_6 ;
wire \top/processor/sha_core/n10755_5 ;
wire \top/processor/sha_core/n10755_6 ;
wire \top/processor/sha_core/n10754_5 ;
wire \top/processor/sha_core/n10754_6 ;
wire \top/processor/sha_core/n10753_5 ;
wire \top/processor/sha_core/n10753_6 ;
wire \top/processor/sha_core/n10752_5 ;
wire \top/processor/sha_core/n10752_1_COUT ;
wire \top/processor/sha_core/n10783_7 ;
wire \top/processor/sha_core/n10783_8 ;
wire \top/processor/sha_core/n10782_7 ;
wire \top/processor/sha_core/n10782_8 ;
wire \top/processor/sha_core/n10781_7 ;
wire \top/processor/sha_core/n10781_8 ;
wire \top/processor/sha_core/n10780_7 ;
wire \top/processor/sha_core/n10780_8 ;
wire \top/processor/sha_core/n10779_7 ;
wire \top/processor/sha_core/n10779_8 ;
wire \top/processor/sha_core/n10778_7 ;
wire \top/processor/sha_core/n10778_8 ;
wire \top/processor/sha_core/n10777_7 ;
wire \top/processor/sha_core/n10777_8 ;
wire \top/processor/sha_core/n10776_7 ;
wire \top/processor/sha_core/n10776_8 ;
wire \top/processor/sha_core/n10775_7 ;
wire \top/processor/sha_core/n10775_8 ;
wire \top/processor/sha_core/n10774_7 ;
wire \top/processor/sha_core/n10774_8 ;
wire \top/processor/sha_core/n10773_7 ;
wire \top/processor/sha_core/n10773_8 ;
wire \top/processor/sha_core/n10772_7 ;
wire \top/processor/sha_core/n10772_8 ;
wire \top/processor/sha_core/n10771_7 ;
wire \top/processor/sha_core/n10771_8 ;
wire \top/processor/sha_core/n10770_7 ;
wire \top/processor/sha_core/n10770_8 ;
wire \top/processor/sha_core/n10769_7 ;
wire \top/processor/sha_core/n10769_8 ;
wire \top/processor/sha_core/n10768_7 ;
wire \top/processor/sha_core/n10768_8 ;
wire \top/processor/sha_core/n10767_7 ;
wire \top/processor/sha_core/n10767_8 ;
wire \top/processor/sha_core/n10766_7 ;
wire \top/processor/sha_core/n10766_8 ;
wire \top/processor/sha_core/n10765_7 ;
wire \top/processor/sha_core/n10765_8 ;
wire \top/processor/sha_core/n10764_7 ;
wire \top/processor/sha_core/n10764_8 ;
wire \top/processor/sha_core/n10763_7 ;
wire \top/processor/sha_core/n10763_8 ;
wire \top/processor/sha_core/n10762_7 ;
wire \top/processor/sha_core/n10762_8 ;
wire \top/processor/sha_core/n10761_7 ;
wire \top/processor/sha_core/n10761_8 ;
wire \top/processor/sha_core/n10760_7 ;
wire \top/processor/sha_core/n10760_8 ;
wire \top/processor/sha_core/n10759_7 ;
wire \top/processor/sha_core/n10759_8 ;
wire \top/processor/sha_core/n10758_7 ;
wire \top/processor/sha_core/n10758_8 ;
wire \top/processor/sha_core/n10757_7 ;
wire \top/processor/sha_core/n10757_8 ;
wire \top/processor/sha_core/n10756_7 ;
wire \top/processor/sha_core/n10756_8 ;
wire \top/processor/sha_core/n10755_7 ;
wire \top/processor/sha_core/n10755_8 ;
wire \top/processor/sha_core/n10754_7 ;
wire \top/processor/sha_core/n10754_8 ;
wire \top/processor/sha_core/n10753_7 ;
wire \top/processor/sha_core/n10753_8 ;
wire \top/processor/sha_core/n10752_7 ;
wire \top/processor/sha_core/n10752_2_COUT ;
wire \top/processor/sha_core/n10783_9 ;
wire \top/processor/sha_core/n10783_10 ;
wire \top/processor/sha_core/n10782_9 ;
wire \top/processor/sha_core/n10782_10 ;
wire \top/processor/sha_core/n10781_9 ;
wire \top/processor/sha_core/n10781_10 ;
wire \top/processor/sha_core/n10780_9 ;
wire \top/processor/sha_core/n10780_10 ;
wire \top/processor/sha_core/n10779_9 ;
wire \top/processor/sha_core/n10779_10 ;
wire \top/processor/sha_core/n10778_9 ;
wire \top/processor/sha_core/n10778_10 ;
wire \top/processor/sha_core/n10777_9 ;
wire \top/processor/sha_core/n10777_10 ;
wire \top/processor/sha_core/n10776_9 ;
wire \top/processor/sha_core/n10776_10 ;
wire \top/processor/sha_core/n10775_9 ;
wire \top/processor/sha_core/n10775_10 ;
wire \top/processor/sha_core/n10774_9 ;
wire \top/processor/sha_core/n10774_10 ;
wire \top/processor/sha_core/n10773_9 ;
wire \top/processor/sha_core/n10773_10 ;
wire \top/processor/sha_core/n10772_9 ;
wire \top/processor/sha_core/n10772_10 ;
wire \top/processor/sha_core/n10771_9 ;
wire \top/processor/sha_core/n10771_10 ;
wire \top/processor/sha_core/n10770_9 ;
wire \top/processor/sha_core/n10770_10 ;
wire \top/processor/sha_core/n10769_9 ;
wire \top/processor/sha_core/n10769_10 ;
wire \top/processor/sha_core/n10768_9 ;
wire \top/processor/sha_core/n10768_10 ;
wire \top/processor/sha_core/n10767_9 ;
wire \top/processor/sha_core/n10767_10 ;
wire \top/processor/sha_core/n10766_9 ;
wire \top/processor/sha_core/n10766_10 ;
wire \top/processor/sha_core/n10765_9 ;
wire \top/processor/sha_core/n10765_10 ;
wire \top/processor/sha_core/n10764_9 ;
wire \top/processor/sha_core/n10764_10 ;
wire \top/processor/sha_core/n10763_9 ;
wire \top/processor/sha_core/n10763_10 ;
wire \top/processor/sha_core/n10762_9 ;
wire \top/processor/sha_core/n10762_10 ;
wire \top/processor/sha_core/n10761_9 ;
wire \top/processor/sha_core/n10761_10 ;
wire \top/processor/sha_core/n10760_9 ;
wire \top/processor/sha_core/n10760_10 ;
wire \top/processor/sha_core/n10759_9 ;
wire \top/processor/sha_core/n10759_10 ;
wire \top/processor/sha_core/n10758_9 ;
wire \top/processor/sha_core/n10758_10 ;
wire \top/processor/sha_core/n10757_9 ;
wire \top/processor/sha_core/n10757_10 ;
wire \top/processor/sha_core/n10756_9 ;
wire \top/processor/sha_core/n10756_10 ;
wire \top/processor/sha_core/n10755_9 ;
wire \top/processor/sha_core/n10755_10 ;
wire \top/processor/sha_core/n10754_9 ;
wire \top/processor/sha_core/n10754_10 ;
wire \top/processor/sha_core/n10753_9 ;
wire \top/processor/sha_core/n10753_10 ;
wire \top/processor/sha_core/n10752_9 ;
wire \top/processor/sha_core/n10752_3_COUT ;
wire \top/processor/sha_core/n10783_11 ;
wire \top/processor/sha_core/n10783_12 ;
wire \top/processor/sha_core/n10782_11 ;
wire \top/processor/sha_core/n10782_12 ;
wire \top/processor/sha_core/n10781_11 ;
wire \top/processor/sha_core/n10781_12 ;
wire \top/processor/sha_core/n10780_11 ;
wire \top/processor/sha_core/n10780_12 ;
wire \top/processor/sha_core/n10779_11 ;
wire \top/processor/sha_core/n10779_12 ;
wire \top/processor/sha_core/n10778_11 ;
wire \top/processor/sha_core/n10778_12 ;
wire \top/processor/sha_core/n10777_11 ;
wire \top/processor/sha_core/n10777_12 ;
wire \top/processor/sha_core/n10776_11 ;
wire \top/processor/sha_core/n10776_12 ;
wire \top/processor/sha_core/n10775_11 ;
wire \top/processor/sha_core/n10775_12 ;
wire \top/processor/sha_core/n10774_11 ;
wire \top/processor/sha_core/n10774_12 ;
wire \top/processor/sha_core/n10773_11 ;
wire \top/processor/sha_core/n10773_12 ;
wire \top/processor/sha_core/n10772_11 ;
wire \top/processor/sha_core/n10772_12 ;
wire \top/processor/sha_core/n10771_11 ;
wire \top/processor/sha_core/n10771_12 ;
wire \top/processor/sha_core/n10770_11 ;
wire \top/processor/sha_core/n10770_12 ;
wire \top/processor/sha_core/n10769_11 ;
wire \top/processor/sha_core/n10769_12 ;
wire \top/processor/sha_core/n10768_11 ;
wire \top/processor/sha_core/n10768_12 ;
wire \top/processor/sha_core/n10767_11 ;
wire \top/processor/sha_core/n10767_12 ;
wire \top/processor/sha_core/n10766_11 ;
wire \top/processor/sha_core/n10766_12 ;
wire \top/processor/sha_core/n10765_11 ;
wire \top/processor/sha_core/n10765_12 ;
wire \top/processor/sha_core/n10764_11 ;
wire \top/processor/sha_core/n10764_12 ;
wire \top/processor/sha_core/n10763_11 ;
wire \top/processor/sha_core/n10763_12 ;
wire \top/processor/sha_core/n10762_11 ;
wire \top/processor/sha_core/n10762_12 ;
wire \top/processor/sha_core/n10761_11 ;
wire \top/processor/sha_core/n10761_12 ;
wire \top/processor/sha_core/n10760_11 ;
wire \top/processor/sha_core/n10760_12 ;
wire \top/processor/sha_core/n10759_11 ;
wire \top/processor/sha_core/n10759_12 ;
wire \top/processor/sha_core/n10758_11 ;
wire \top/processor/sha_core/n10758_12 ;
wire \top/processor/sha_core/n10757_11 ;
wire \top/processor/sha_core/n10757_12 ;
wire \top/processor/sha_core/n10756_11 ;
wire \top/processor/sha_core/n10756_12 ;
wire \top/processor/sha_core/n10755_11 ;
wire \top/processor/sha_core/n10755_12 ;
wire \top/processor/sha_core/n10754_11 ;
wire \top/processor/sha_core/n10754_12 ;
wire \top/processor/sha_core/n10753_11 ;
wire \top/processor/sha_core/n10753_12 ;
wire \top/processor/sha_core/n10752_11 ;
wire \top/processor/sha_core/n10752_4_COUT ;
wire \top/processor/sha_core/n10816_3 ;
wire \top/processor/sha_core/n10816_4 ;
wire \top/processor/sha_core/n10815_3 ;
wire \top/processor/sha_core/n10815_4 ;
wire \top/processor/sha_core/n10814_3 ;
wire \top/processor/sha_core/n10814_4 ;
wire \top/processor/sha_core/n10813_3 ;
wire \top/processor/sha_core/n10813_4 ;
wire \top/processor/sha_core/n10812_3 ;
wire \top/processor/sha_core/n10812_4 ;
wire \top/processor/sha_core/n10811_3 ;
wire \top/processor/sha_core/n10811_4 ;
wire \top/processor/sha_core/n10810_3 ;
wire \top/processor/sha_core/n10810_4 ;
wire \top/processor/sha_core/n10809_3 ;
wire \top/processor/sha_core/n10809_4 ;
wire \top/processor/sha_core/n10808_3 ;
wire \top/processor/sha_core/n10808_4 ;
wire \top/processor/sha_core/n10807_3 ;
wire \top/processor/sha_core/n10807_4 ;
wire \top/processor/sha_core/n10806_3 ;
wire \top/processor/sha_core/n10806_4 ;
wire \top/processor/sha_core/n10805_3 ;
wire \top/processor/sha_core/n10805_4 ;
wire \top/processor/sha_core/n10804_3 ;
wire \top/processor/sha_core/n10804_4 ;
wire \top/processor/sha_core/n10803_3 ;
wire \top/processor/sha_core/n10803_4 ;
wire \top/processor/sha_core/n10802_3 ;
wire \top/processor/sha_core/n10802_4 ;
wire \top/processor/sha_core/n10801_3 ;
wire \top/processor/sha_core/n10801_4 ;
wire \top/processor/sha_core/n10800_3 ;
wire \top/processor/sha_core/n10800_4 ;
wire \top/processor/sha_core/n10799_3 ;
wire \top/processor/sha_core/n10799_4 ;
wire \top/processor/sha_core/n10798_3 ;
wire \top/processor/sha_core/n10798_4 ;
wire \top/processor/sha_core/n10797_3 ;
wire \top/processor/sha_core/n10797_4 ;
wire \top/processor/sha_core/n10796_3 ;
wire \top/processor/sha_core/n10796_4 ;
wire \top/processor/sha_core/n10795_3 ;
wire \top/processor/sha_core/n10795_4 ;
wire \top/processor/sha_core/n10794_3 ;
wire \top/processor/sha_core/n10794_4 ;
wire \top/processor/sha_core/n10793_3 ;
wire \top/processor/sha_core/n10793_4 ;
wire \top/processor/sha_core/n10792_3 ;
wire \top/processor/sha_core/n10792_4 ;
wire \top/processor/sha_core/n10791_3 ;
wire \top/processor/sha_core/n10791_4 ;
wire \top/processor/sha_core/n10790_3 ;
wire \top/processor/sha_core/n10790_4 ;
wire \top/processor/sha_core/n10789_3 ;
wire \top/processor/sha_core/n10789_4 ;
wire \top/processor/sha_core/n10788_3 ;
wire \top/processor/sha_core/n10788_4 ;
wire \top/processor/sha_core/n10787_3 ;
wire \top/processor/sha_core/n10787_4 ;
wire \top/processor/sha_core/n10786_3 ;
wire \top/processor/sha_core/n10786_4 ;
wire \top/processor/sha_core/n10785_3 ;
wire \top/processor/sha_core/n10785_0_COUT ;
wire \top/processor/sha_core/n10816_5 ;
wire \top/processor/sha_core/n10816_6 ;
wire \top/processor/sha_core/n10815_5 ;
wire \top/processor/sha_core/n10815_6 ;
wire \top/processor/sha_core/n10814_5 ;
wire \top/processor/sha_core/n10814_6 ;
wire \top/processor/sha_core/n10813_5 ;
wire \top/processor/sha_core/n10813_6 ;
wire \top/processor/sha_core/n10812_5 ;
wire \top/processor/sha_core/n10812_6 ;
wire \top/processor/sha_core/n10811_5 ;
wire \top/processor/sha_core/n10811_6 ;
wire \top/processor/sha_core/n10810_5 ;
wire \top/processor/sha_core/n10810_6 ;
wire \top/processor/sha_core/n10809_5 ;
wire \top/processor/sha_core/n10809_6 ;
wire \top/processor/sha_core/n10808_5 ;
wire \top/processor/sha_core/n10808_6 ;
wire \top/processor/sha_core/n10807_5 ;
wire \top/processor/sha_core/n10807_6 ;
wire \top/processor/sha_core/n10806_5 ;
wire \top/processor/sha_core/n10806_6 ;
wire \top/processor/sha_core/n10805_5 ;
wire \top/processor/sha_core/n10805_6 ;
wire \top/processor/sha_core/n10804_5 ;
wire \top/processor/sha_core/n10804_6 ;
wire \top/processor/sha_core/n10803_5 ;
wire \top/processor/sha_core/n10803_6 ;
wire \top/processor/sha_core/n10802_5 ;
wire \top/processor/sha_core/n10802_6 ;
wire \top/processor/sha_core/n10801_5 ;
wire \top/processor/sha_core/n10801_6 ;
wire \top/processor/sha_core/n10800_5 ;
wire \top/processor/sha_core/n10800_6 ;
wire \top/processor/sha_core/n10799_5 ;
wire \top/processor/sha_core/n10799_6 ;
wire \top/processor/sha_core/n10798_5 ;
wire \top/processor/sha_core/n10798_6 ;
wire \top/processor/sha_core/n10797_5 ;
wire \top/processor/sha_core/n10797_6 ;
wire \top/processor/sha_core/n10796_5 ;
wire \top/processor/sha_core/n10796_6 ;
wire \top/processor/sha_core/n10795_5 ;
wire \top/processor/sha_core/n10795_6 ;
wire \top/processor/sha_core/n10794_5 ;
wire \top/processor/sha_core/n10794_6 ;
wire \top/processor/sha_core/n10793_5 ;
wire \top/processor/sha_core/n10793_6 ;
wire \top/processor/sha_core/n10792_5 ;
wire \top/processor/sha_core/n10792_6 ;
wire \top/processor/sha_core/n10791_5 ;
wire \top/processor/sha_core/n10791_6 ;
wire \top/processor/sha_core/n10790_5 ;
wire \top/processor/sha_core/n10790_6 ;
wire \top/processor/sha_core/n10789_5 ;
wire \top/processor/sha_core/n10789_6 ;
wire \top/processor/sha_core/n10788_5 ;
wire \top/processor/sha_core/n10788_6 ;
wire \top/processor/sha_core/n10787_5 ;
wire \top/processor/sha_core/n10787_6 ;
wire \top/processor/sha_core/n10786_5 ;
wire \top/processor/sha_core/n10786_6 ;
wire \top/processor/sha_core/n10785_5 ;
wire \top/processor/sha_core/n10785_1_COUT ;
wire \top/processor/sha_core/n10816_7 ;
wire \top/processor/sha_core/n10816_8 ;
wire \top/processor/sha_core/n10815_7 ;
wire \top/processor/sha_core/n10815_8 ;
wire \top/processor/sha_core/n10814_7 ;
wire \top/processor/sha_core/n10814_8 ;
wire \top/processor/sha_core/n10813_7 ;
wire \top/processor/sha_core/n10813_8 ;
wire \top/processor/sha_core/n10812_7 ;
wire \top/processor/sha_core/n10812_8 ;
wire \top/processor/sha_core/n10811_7 ;
wire \top/processor/sha_core/n10811_8 ;
wire \top/processor/sha_core/n10810_7 ;
wire \top/processor/sha_core/n10810_8 ;
wire \top/processor/sha_core/n10809_7 ;
wire \top/processor/sha_core/n10809_8 ;
wire \top/processor/sha_core/n10808_7 ;
wire \top/processor/sha_core/n10808_8 ;
wire \top/processor/sha_core/n10807_7 ;
wire \top/processor/sha_core/n10807_8 ;
wire \top/processor/sha_core/n10806_7 ;
wire \top/processor/sha_core/n10806_8 ;
wire \top/processor/sha_core/n10805_7 ;
wire \top/processor/sha_core/n10805_8 ;
wire \top/processor/sha_core/n10804_7 ;
wire \top/processor/sha_core/n10804_8 ;
wire \top/processor/sha_core/n10803_7 ;
wire \top/processor/sha_core/n10803_8 ;
wire \top/processor/sha_core/n10802_7 ;
wire \top/processor/sha_core/n10802_8 ;
wire \top/processor/sha_core/n10801_7 ;
wire \top/processor/sha_core/n10801_8 ;
wire \top/processor/sha_core/n10800_7 ;
wire \top/processor/sha_core/n10800_8 ;
wire \top/processor/sha_core/n10799_7 ;
wire \top/processor/sha_core/n10799_8 ;
wire \top/processor/sha_core/n10798_7 ;
wire \top/processor/sha_core/n10798_8 ;
wire \top/processor/sha_core/n10797_7 ;
wire \top/processor/sha_core/n10797_8 ;
wire \top/processor/sha_core/n10796_7 ;
wire \top/processor/sha_core/n10796_8 ;
wire \top/processor/sha_core/n10795_7 ;
wire \top/processor/sha_core/n10795_8 ;
wire \top/processor/sha_core/n10794_7 ;
wire \top/processor/sha_core/n10794_8 ;
wire \top/processor/sha_core/n10793_7 ;
wire \top/processor/sha_core/n10793_8 ;
wire \top/processor/sha_core/n10792_7 ;
wire \top/processor/sha_core/n10792_8 ;
wire \top/processor/sha_core/n10791_7 ;
wire \top/processor/sha_core/n10791_8 ;
wire \top/processor/sha_core/n10790_7 ;
wire \top/processor/sha_core/n10790_8 ;
wire \top/processor/sha_core/n10789_7 ;
wire \top/processor/sha_core/n10789_8 ;
wire \top/processor/sha_core/n10788_7 ;
wire \top/processor/sha_core/n10788_8 ;
wire \top/processor/sha_core/n10787_7 ;
wire \top/processor/sha_core/n10787_8 ;
wire \top/processor/sha_core/n10786_7 ;
wire \top/processor/sha_core/n10786_8 ;
wire \top/processor/sha_core/n10785_7 ;
wire \top/processor/sha_core/n10785_2_COUT ;
wire \top/processor/sha_core/n10816_9 ;
wire \top/processor/sha_core/n10816_10 ;
wire \top/processor/sha_core/n10815_9 ;
wire \top/processor/sha_core/n10815_10 ;
wire \top/processor/sha_core/n10814_9 ;
wire \top/processor/sha_core/n10814_10 ;
wire \top/processor/sha_core/n10813_9 ;
wire \top/processor/sha_core/n10813_10 ;
wire \top/processor/sha_core/n10812_9 ;
wire \top/processor/sha_core/n10812_10 ;
wire \top/processor/sha_core/n10811_9 ;
wire \top/processor/sha_core/n10811_10 ;
wire \top/processor/sha_core/n10810_9 ;
wire \top/processor/sha_core/n10810_10 ;
wire \top/processor/sha_core/n10809_9 ;
wire \top/processor/sha_core/n10809_10 ;
wire \top/processor/sha_core/n10808_9 ;
wire \top/processor/sha_core/n10808_10 ;
wire \top/processor/sha_core/n10807_9 ;
wire \top/processor/sha_core/n10807_10 ;
wire \top/processor/sha_core/n10806_9 ;
wire \top/processor/sha_core/n10806_10 ;
wire \top/processor/sha_core/n10805_9 ;
wire \top/processor/sha_core/n10805_10 ;
wire \top/processor/sha_core/n10804_9 ;
wire \top/processor/sha_core/n10804_10 ;
wire \top/processor/sha_core/n10803_9 ;
wire \top/processor/sha_core/n10803_10 ;
wire \top/processor/sha_core/n10802_9 ;
wire \top/processor/sha_core/n10802_10 ;
wire \top/processor/sha_core/n10801_9 ;
wire \top/processor/sha_core/n10801_10 ;
wire \top/processor/sha_core/n10800_9 ;
wire \top/processor/sha_core/n10800_10 ;
wire \top/processor/sha_core/n10799_9 ;
wire \top/processor/sha_core/n10799_10 ;
wire \top/processor/sha_core/n10798_9 ;
wire \top/processor/sha_core/n10798_10 ;
wire \top/processor/sha_core/n10797_9 ;
wire \top/processor/sha_core/n10797_10 ;
wire \top/processor/sha_core/n10796_9 ;
wire \top/processor/sha_core/n10796_10 ;
wire \top/processor/sha_core/n10795_9 ;
wire \top/processor/sha_core/n10795_10 ;
wire \top/processor/sha_core/n10794_9 ;
wire \top/processor/sha_core/n10794_10 ;
wire \top/processor/sha_core/n10793_9 ;
wire \top/processor/sha_core/n10793_10 ;
wire \top/processor/sha_core/n10792_9 ;
wire \top/processor/sha_core/n10792_10 ;
wire \top/processor/sha_core/n10791_9 ;
wire \top/processor/sha_core/n10791_10 ;
wire \top/processor/sha_core/n10790_9 ;
wire \top/processor/sha_core/n10790_10 ;
wire \top/processor/sha_core/n10789_9 ;
wire \top/processor/sha_core/n10789_10 ;
wire \top/processor/sha_core/n10788_9 ;
wire \top/processor/sha_core/n10788_10 ;
wire \top/processor/sha_core/n10787_9 ;
wire \top/processor/sha_core/n10787_10 ;
wire \top/processor/sha_core/n10786_9 ;
wire \top/processor/sha_core/n10786_10 ;
wire \top/processor/sha_core/n10785_9 ;
wire \top/processor/sha_core/n10785_3_COUT ;
wire \top/processor/sha_core/n10816_11 ;
wire \top/processor/sha_core/n10816_12 ;
wire \top/processor/sha_core/n10815_11 ;
wire \top/processor/sha_core/n10815_12 ;
wire \top/processor/sha_core/n10814_11 ;
wire \top/processor/sha_core/n10814_12 ;
wire \top/processor/sha_core/n10813_11 ;
wire \top/processor/sha_core/n10813_12 ;
wire \top/processor/sha_core/n10812_11 ;
wire \top/processor/sha_core/n10812_12 ;
wire \top/processor/sha_core/n10811_11 ;
wire \top/processor/sha_core/n10811_12 ;
wire \top/processor/sha_core/n10810_11 ;
wire \top/processor/sha_core/n10810_12 ;
wire \top/processor/sha_core/n10809_11 ;
wire \top/processor/sha_core/n10809_12 ;
wire \top/processor/sha_core/n10808_11 ;
wire \top/processor/sha_core/n10808_12 ;
wire \top/processor/sha_core/n10807_11 ;
wire \top/processor/sha_core/n10807_12 ;
wire \top/processor/sha_core/n10806_11 ;
wire \top/processor/sha_core/n10806_12 ;
wire \top/processor/sha_core/n10805_11 ;
wire \top/processor/sha_core/n10805_12 ;
wire \top/processor/sha_core/n10804_11 ;
wire \top/processor/sha_core/n10804_12 ;
wire \top/processor/sha_core/n10803_11 ;
wire \top/processor/sha_core/n10803_12 ;
wire \top/processor/sha_core/n10802_11 ;
wire \top/processor/sha_core/n10802_12 ;
wire \top/processor/sha_core/n10801_11 ;
wire \top/processor/sha_core/n10801_12 ;
wire \top/processor/sha_core/n10800_11 ;
wire \top/processor/sha_core/n10800_12 ;
wire \top/processor/sha_core/n10799_11 ;
wire \top/processor/sha_core/n10799_12 ;
wire \top/processor/sha_core/n10798_11 ;
wire \top/processor/sha_core/n10798_12 ;
wire \top/processor/sha_core/n10797_11 ;
wire \top/processor/sha_core/n10797_12 ;
wire \top/processor/sha_core/n10796_11 ;
wire \top/processor/sha_core/n10796_12 ;
wire \top/processor/sha_core/n10795_11 ;
wire \top/processor/sha_core/n10795_12 ;
wire \top/processor/sha_core/n10794_11 ;
wire \top/processor/sha_core/n10794_12 ;
wire \top/processor/sha_core/n10793_11 ;
wire \top/processor/sha_core/n10793_12 ;
wire \top/processor/sha_core/n10792_11 ;
wire \top/processor/sha_core/n10792_12 ;
wire \top/processor/sha_core/n10791_11 ;
wire \top/processor/sha_core/n10791_12 ;
wire \top/processor/sha_core/n10790_11 ;
wire \top/processor/sha_core/n10790_12 ;
wire \top/processor/sha_core/n10789_11 ;
wire \top/processor/sha_core/n10789_12 ;
wire \top/processor/sha_core/n10788_11 ;
wire \top/processor/sha_core/n10788_12 ;
wire \top/processor/sha_core/n10787_11 ;
wire \top/processor/sha_core/n10787_12 ;
wire \top/processor/sha_core/n10786_11 ;
wire \top/processor/sha_core/n10786_12 ;
wire \top/processor/sha_core/n10785_11 ;
wire \top/processor/sha_core/n10785_4_COUT ;
wire \top/processor/sha_core/n10816_13 ;
wire \top/processor/sha_core/n10816_14 ;
wire \top/processor/sha_core/n10815_13 ;
wire \top/processor/sha_core/n10815_14 ;
wire \top/processor/sha_core/n10814_13 ;
wire \top/processor/sha_core/n10814_14 ;
wire \top/processor/sha_core/n10813_13 ;
wire \top/processor/sha_core/n10813_14 ;
wire \top/processor/sha_core/n10812_13 ;
wire \top/processor/sha_core/n10812_14 ;
wire \top/processor/sha_core/n10811_13 ;
wire \top/processor/sha_core/n10811_14 ;
wire \top/processor/sha_core/n10810_13 ;
wire \top/processor/sha_core/n10810_14 ;
wire \top/processor/sha_core/n10809_13 ;
wire \top/processor/sha_core/n10809_14 ;
wire \top/processor/sha_core/n10808_13 ;
wire \top/processor/sha_core/n10808_14 ;
wire \top/processor/sha_core/n10807_13 ;
wire \top/processor/sha_core/n10807_14 ;
wire \top/processor/sha_core/n10806_13 ;
wire \top/processor/sha_core/n10806_14 ;
wire \top/processor/sha_core/n10805_13 ;
wire \top/processor/sha_core/n10805_14 ;
wire \top/processor/sha_core/n10804_13 ;
wire \top/processor/sha_core/n10804_14 ;
wire \top/processor/sha_core/n10803_13 ;
wire \top/processor/sha_core/n10803_14 ;
wire \top/processor/sha_core/n10802_13 ;
wire \top/processor/sha_core/n10802_14 ;
wire \top/processor/sha_core/n10801_13 ;
wire \top/processor/sha_core/n10801_14 ;
wire \top/processor/sha_core/n10800_13 ;
wire \top/processor/sha_core/n10800_14 ;
wire \top/processor/sha_core/n10799_13 ;
wire \top/processor/sha_core/n10799_14 ;
wire \top/processor/sha_core/n10798_13 ;
wire \top/processor/sha_core/n10798_14 ;
wire \top/processor/sha_core/n10797_13 ;
wire \top/processor/sha_core/n10797_14 ;
wire \top/processor/sha_core/n10796_13 ;
wire \top/processor/sha_core/n10796_14 ;
wire \top/processor/sha_core/n10795_13 ;
wire \top/processor/sha_core/n10795_14 ;
wire \top/processor/sha_core/n10794_13 ;
wire \top/processor/sha_core/n10794_14 ;
wire \top/processor/sha_core/n10793_13 ;
wire \top/processor/sha_core/n10793_14 ;
wire \top/processor/sha_core/n10792_13 ;
wire \top/processor/sha_core/n10792_14 ;
wire \top/processor/sha_core/n10791_13 ;
wire \top/processor/sha_core/n10791_14 ;
wire \top/processor/sha_core/n10790_13 ;
wire \top/processor/sha_core/n10790_14 ;
wire \top/processor/sha_core/n10789_13 ;
wire \top/processor/sha_core/n10789_14 ;
wire \top/processor/sha_core/n10788_13 ;
wire \top/processor/sha_core/n10788_14 ;
wire \top/processor/sha_core/n10787_13 ;
wire \top/processor/sha_core/n10787_14 ;
wire \top/processor/sha_core/n10786_13 ;
wire \top/processor/sha_core/n10786_14 ;
wire \top/processor/sha_core/n10785_13 ;
wire \top/processor/sha_core/n10785_5_COUT ;
wire \top/processor/sha_core/n327_165 ;
wire \top/processor/sha_core/n327_167 ;
wire \top/processor/sha_core/n327_169 ;
wire \top/processor/sha_core/n327_171 ;
wire \top/processor/sha_core/n327_173 ;
wire \top/processor/sha_core/n327_175 ;
wire \top/processor/sha_core/n327_177 ;
wire \top/processor/sha_core/n327_179 ;
wire \top/processor/sha_core/n327_181 ;
wire \top/processor/sha_core/n327_183 ;
wire \top/processor/sha_core/n327_185 ;
wire \top/processor/sha_core/n327_187 ;
wire \top/processor/sha_core/n327_189 ;
wire \top/processor/sha_core/n327_191 ;
wire \top/processor/sha_core/n327_193 ;
wire \top/processor/sha_core/n327_195 ;
wire \top/processor/sha_core/n328_165 ;
wire \top/processor/sha_core/n328_167 ;
wire \top/processor/sha_core/n328_169 ;
wire \top/processor/sha_core/n328_171 ;
wire \top/processor/sha_core/n328_173 ;
wire \top/processor/sha_core/n328_175 ;
wire \top/processor/sha_core/n328_177 ;
wire \top/processor/sha_core/n328_179 ;
wire \top/processor/sha_core/n328_181 ;
wire \top/processor/sha_core/n328_183 ;
wire \top/processor/sha_core/n328_185 ;
wire \top/processor/sha_core/n328_187 ;
wire \top/processor/sha_core/n328_189 ;
wire \top/processor/sha_core/n328_191 ;
wire \top/processor/sha_core/n328_193 ;
wire \top/processor/sha_core/n328_195 ;
wire \top/processor/sha_core/n329_165 ;
wire \top/processor/sha_core/n329_167 ;
wire \top/processor/sha_core/n329_169 ;
wire \top/processor/sha_core/n329_171 ;
wire \top/processor/sha_core/n329_173 ;
wire \top/processor/sha_core/n329_175 ;
wire \top/processor/sha_core/n329_177 ;
wire \top/processor/sha_core/n329_179 ;
wire \top/processor/sha_core/n329_181 ;
wire \top/processor/sha_core/n329_183 ;
wire \top/processor/sha_core/n329_185 ;
wire \top/processor/sha_core/n329_187 ;
wire \top/processor/sha_core/n329_189 ;
wire \top/processor/sha_core/n329_191 ;
wire \top/processor/sha_core/n329_193 ;
wire \top/processor/sha_core/n329_195 ;
wire \top/processor/sha_core/n330_165 ;
wire \top/processor/sha_core/n330_167 ;
wire \top/processor/sha_core/n330_169 ;
wire \top/processor/sha_core/n330_171 ;
wire \top/processor/sha_core/n330_173 ;
wire \top/processor/sha_core/n330_175 ;
wire \top/processor/sha_core/n330_177 ;
wire \top/processor/sha_core/n330_179 ;
wire \top/processor/sha_core/n330_181 ;
wire \top/processor/sha_core/n330_183 ;
wire \top/processor/sha_core/n330_185 ;
wire \top/processor/sha_core/n330_187 ;
wire \top/processor/sha_core/n330_189 ;
wire \top/processor/sha_core/n330_191 ;
wire \top/processor/sha_core/n330_193 ;
wire \top/processor/sha_core/n330_195 ;
wire \top/processor/sha_core/n331_165 ;
wire \top/processor/sha_core/n331_167 ;
wire \top/processor/sha_core/n331_169 ;
wire \top/processor/sha_core/n331_171 ;
wire \top/processor/sha_core/n331_173 ;
wire \top/processor/sha_core/n331_175 ;
wire \top/processor/sha_core/n331_177 ;
wire \top/processor/sha_core/n331_179 ;
wire \top/processor/sha_core/n331_181 ;
wire \top/processor/sha_core/n331_183 ;
wire \top/processor/sha_core/n331_185 ;
wire \top/processor/sha_core/n331_187 ;
wire \top/processor/sha_core/n331_189 ;
wire \top/processor/sha_core/n331_191 ;
wire \top/processor/sha_core/n331_193 ;
wire \top/processor/sha_core/n331_195 ;
wire \top/processor/sha_core/n332_165 ;
wire \top/processor/sha_core/n332_167 ;
wire \top/processor/sha_core/n332_169 ;
wire \top/processor/sha_core/n332_171 ;
wire \top/processor/sha_core/n332_173 ;
wire \top/processor/sha_core/n332_175 ;
wire \top/processor/sha_core/n332_177 ;
wire \top/processor/sha_core/n332_179 ;
wire \top/processor/sha_core/n332_181 ;
wire \top/processor/sha_core/n332_183 ;
wire \top/processor/sha_core/n332_185 ;
wire \top/processor/sha_core/n332_187 ;
wire \top/processor/sha_core/n332_189 ;
wire \top/processor/sha_core/n332_191 ;
wire \top/processor/sha_core/n332_193 ;
wire \top/processor/sha_core/n332_195 ;
wire \top/processor/sha_core/n333_165 ;
wire \top/processor/sha_core/n333_167 ;
wire \top/processor/sha_core/n333_169 ;
wire \top/processor/sha_core/n333_171 ;
wire \top/processor/sha_core/n333_173 ;
wire \top/processor/sha_core/n333_175 ;
wire \top/processor/sha_core/n333_177 ;
wire \top/processor/sha_core/n333_179 ;
wire \top/processor/sha_core/n333_181 ;
wire \top/processor/sha_core/n333_183 ;
wire \top/processor/sha_core/n333_185 ;
wire \top/processor/sha_core/n333_187 ;
wire \top/processor/sha_core/n333_189 ;
wire \top/processor/sha_core/n333_191 ;
wire \top/processor/sha_core/n333_193 ;
wire \top/processor/sha_core/n333_195 ;
wire \top/processor/sha_core/n334_165 ;
wire \top/processor/sha_core/n334_167 ;
wire \top/processor/sha_core/n334_169 ;
wire \top/processor/sha_core/n334_171 ;
wire \top/processor/sha_core/n334_173 ;
wire \top/processor/sha_core/n334_175 ;
wire \top/processor/sha_core/n334_177 ;
wire \top/processor/sha_core/n334_179 ;
wire \top/processor/sha_core/n334_181 ;
wire \top/processor/sha_core/n334_183 ;
wire \top/processor/sha_core/n334_185 ;
wire \top/processor/sha_core/n334_187 ;
wire \top/processor/sha_core/n334_189 ;
wire \top/processor/sha_core/n334_191 ;
wire \top/processor/sha_core/n334_193 ;
wire \top/processor/sha_core/n334_195 ;
wire \top/processor/sha_core/n335_165 ;
wire \top/processor/sha_core/n335_167 ;
wire \top/processor/sha_core/n335_169 ;
wire \top/processor/sha_core/n335_171 ;
wire \top/processor/sha_core/n335_173 ;
wire \top/processor/sha_core/n335_175 ;
wire \top/processor/sha_core/n335_177 ;
wire \top/processor/sha_core/n335_179 ;
wire \top/processor/sha_core/n335_181 ;
wire \top/processor/sha_core/n335_183 ;
wire \top/processor/sha_core/n335_185 ;
wire \top/processor/sha_core/n335_187 ;
wire \top/processor/sha_core/n335_189 ;
wire \top/processor/sha_core/n335_191 ;
wire \top/processor/sha_core/n335_193 ;
wire \top/processor/sha_core/n335_195 ;
wire \top/processor/sha_core/n336_165 ;
wire \top/processor/sha_core/n336_167 ;
wire \top/processor/sha_core/n336_169 ;
wire \top/processor/sha_core/n336_171 ;
wire \top/processor/sha_core/n336_173 ;
wire \top/processor/sha_core/n336_175 ;
wire \top/processor/sha_core/n336_177 ;
wire \top/processor/sha_core/n336_179 ;
wire \top/processor/sha_core/n336_181 ;
wire \top/processor/sha_core/n336_183 ;
wire \top/processor/sha_core/n336_185 ;
wire \top/processor/sha_core/n336_187 ;
wire \top/processor/sha_core/n336_189 ;
wire \top/processor/sha_core/n336_191 ;
wire \top/processor/sha_core/n336_193 ;
wire \top/processor/sha_core/n336_195 ;
wire \top/processor/sha_core/n337_165 ;
wire \top/processor/sha_core/n337_167 ;
wire \top/processor/sha_core/n337_169 ;
wire \top/processor/sha_core/n337_171 ;
wire \top/processor/sha_core/n337_173 ;
wire \top/processor/sha_core/n337_175 ;
wire \top/processor/sha_core/n337_177 ;
wire \top/processor/sha_core/n337_179 ;
wire \top/processor/sha_core/n337_181 ;
wire \top/processor/sha_core/n337_183 ;
wire \top/processor/sha_core/n337_185 ;
wire \top/processor/sha_core/n337_187 ;
wire \top/processor/sha_core/n337_189 ;
wire \top/processor/sha_core/n337_191 ;
wire \top/processor/sha_core/n337_193 ;
wire \top/processor/sha_core/n337_195 ;
wire \top/processor/sha_core/n338_165 ;
wire \top/processor/sha_core/n338_167 ;
wire \top/processor/sha_core/n338_169 ;
wire \top/processor/sha_core/n338_171 ;
wire \top/processor/sha_core/n338_173 ;
wire \top/processor/sha_core/n338_175 ;
wire \top/processor/sha_core/n338_177 ;
wire \top/processor/sha_core/n338_179 ;
wire \top/processor/sha_core/n338_181 ;
wire \top/processor/sha_core/n338_183 ;
wire \top/processor/sha_core/n338_185 ;
wire \top/processor/sha_core/n338_187 ;
wire \top/processor/sha_core/n338_189 ;
wire \top/processor/sha_core/n338_191 ;
wire \top/processor/sha_core/n338_193 ;
wire \top/processor/sha_core/n338_195 ;
wire \top/processor/sha_core/n339_165 ;
wire \top/processor/sha_core/n339_167 ;
wire \top/processor/sha_core/n339_169 ;
wire \top/processor/sha_core/n339_171 ;
wire \top/processor/sha_core/n339_173 ;
wire \top/processor/sha_core/n339_175 ;
wire \top/processor/sha_core/n339_177 ;
wire \top/processor/sha_core/n339_179 ;
wire \top/processor/sha_core/n339_181 ;
wire \top/processor/sha_core/n339_183 ;
wire \top/processor/sha_core/n339_185 ;
wire \top/processor/sha_core/n339_187 ;
wire \top/processor/sha_core/n339_189 ;
wire \top/processor/sha_core/n339_191 ;
wire \top/processor/sha_core/n339_193 ;
wire \top/processor/sha_core/n339_195 ;
wire \top/processor/sha_core/n340_165 ;
wire \top/processor/sha_core/n340_167 ;
wire \top/processor/sha_core/n340_169 ;
wire \top/processor/sha_core/n340_171 ;
wire \top/processor/sha_core/n340_173 ;
wire \top/processor/sha_core/n340_175 ;
wire \top/processor/sha_core/n340_177 ;
wire \top/processor/sha_core/n340_179 ;
wire \top/processor/sha_core/n340_181 ;
wire \top/processor/sha_core/n340_183 ;
wire \top/processor/sha_core/n340_185 ;
wire \top/processor/sha_core/n340_187 ;
wire \top/processor/sha_core/n340_189 ;
wire \top/processor/sha_core/n340_191 ;
wire \top/processor/sha_core/n340_193 ;
wire \top/processor/sha_core/n340_195 ;
wire \top/processor/sha_core/n341_165 ;
wire \top/processor/sha_core/n341_167 ;
wire \top/processor/sha_core/n341_169 ;
wire \top/processor/sha_core/n341_171 ;
wire \top/processor/sha_core/n341_173 ;
wire \top/processor/sha_core/n341_175 ;
wire \top/processor/sha_core/n341_177 ;
wire \top/processor/sha_core/n341_179 ;
wire \top/processor/sha_core/n341_181 ;
wire \top/processor/sha_core/n341_183 ;
wire \top/processor/sha_core/n341_185 ;
wire \top/processor/sha_core/n341_187 ;
wire \top/processor/sha_core/n341_189 ;
wire \top/processor/sha_core/n341_191 ;
wire \top/processor/sha_core/n341_193 ;
wire \top/processor/sha_core/n341_195 ;
wire \top/processor/sha_core/n342_165 ;
wire \top/processor/sha_core/n342_167 ;
wire \top/processor/sha_core/n342_169 ;
wire \top/processor/sha_core/n342_171 ;
wire \top/processor/sha_core/n342_173 ;
wire \top/processor/sha_core/n342_175 ;
wire \top/processor/sha_core/n342_177 ;
wire \top/processor/sha_core/n342_179 ;
wire \top/processor/sha_core/n342_181 ;
wire \top/processor/sha_core/n342_183 ;
wire \top/processor/sha_core/n342_185 ;
wire \top/processor/sha_core/n342_187 ;
wire \top/processor/sha_core/n342_189 ;
wire \top/processor/sha_core/n342_191 ;
wire \top/processor/sha_core/n342_193 ;
wire \top/processor/sha_core/n342_195 ;
wire \top/processor/sha_core/n343_165 ;
wire \top/processor/sha_core/n343_167 ;
wire \top/processor/sha_core/n343_169 ;
wire \top/processor/sha_core/n343_171 ;
wire \top/processor/sha_core/n343_173 ;
wire \top/processor/sha_core/n343_175 ;
wire \top/processor/sha_core/n343_177 ;
wire \top/processor/sha_core/n343_179 ;
wire \top/processor/sha_core/n343_181 ;
wire \top/processor/sha_core/n343_183 ;
wire \top/processor/sha_core/n343_185 ;
wire \top/processor/sha_core/n343_187 ;
wire \top/processor/sha_core/n343_189 ;
wire \top/processor/sha_core/n343_191 ;
wire \top/processor/sha_core/n343_193 ;
wire \top/processor/sha_core/n343_195 ;
wire \top/processor/sha_core/n344_165 ;
wire \top/processor/sha_core/n344_167 ;
wire \top/processor/sha_core/n344_169 ;
wire \top/processor/sha_core/n344_171 ;
wire \top/processor/sha_core/n344_173 ;
wire \top/processor/sha_core/n344_175 ;
wire \top/processor/sha_core/n344_177 ;
wire \top/processor/sha_core/n344_179 ;
wire \top/processor/sha_core/n344_181 ;
wire \top/processor/sha_core/n344_183 ;
wire \top/processor/sha_core/n344_185 ;
wire \top/processor/sha_core/n344_187 ;
wire \top/processor/sha_core/n344_189 ;
wire \top/processor/sha_core/n344_191 ;
wire \top/processor/sha_core/n344_193 ;
wire \top/processor/sha_core/n344_195 ;
wire \top/processor/sha_core/n345_165 ;
wire \top/processor/sha_core/n345_167 ;
wire \top/processor/sha_core/n345_169 ;
wire \top/processor/sha_core/n345_171 ;
wire \top/processor/sha_core/n345_173 ;
wire \top/processor/sha_core/n345_175 ;
wire \top/processor/sha_core/n345_177 ;
wire \top/processor/sha_core/n345_179 ;
wire \top/processor/sha_core/n345_181 ;
wire \top/processor/sha_core/n345_183 ;
wire \top/processor/sha_core/n345_185 ;
wire \top/processor/sha_core/n345_187 ;
wire \top/processor/sha_core/n345_189 ;
wire \top/processor/sha_core/n345_191 ;
wire \top/processor/sha_core/n345_193 ;
wire \top/processor/sha_core/n345_195 ;
wire \top/processor/sha_core/n346_165 ;
wire \top/processor/sha_core/n346_167 ;
wire \top/processor/sha_core/n346_169 ;
wire \top/processor/sha_core/n346_171 ;
wire \top/processor/sha_core/n346_173 ;
wire \top/processor/sha_core/n346_175 ;
wire \top/processor/sha_core/n346_177 ;
wire \top/processor/sha_core/n346_179 ;
wire \top/processor/sha_core/n346_181 ;
wire \top/processor/sha_core/n346_183 ;
wire \top/processor/sha_core/n346_185 ;
wire \top/processor/sha_core/n346_187 ;
wire \top/processor/sha_core/n346_189 ;
wire \top/processor/sha_core/n346_191 ;
wire \top/processor/sha_core/n346_193 ;
wire \top/processor/sha_core/n346_195 ;
wire \top/processor/sha_core/n347_165 ;
wire \top/processor/sha_core/n347_167 ;
wire \top/processor/sha_core/n347_169 ;
wire \top/processor/sha_core/n347_171 ;
wire \top/processor/sha_core/n347_173 ;
wire \top/processor/sha_core/n347_175 ;
wire \top/processor/sha_core/n347_177 ;
wire \top/processor/sha_core/n347_179 ;
wire \top/processor/sha_core/n347_181 ;
wire \top/processor/sha_core/n347_183 ;
wire \top/processor/sha_core/n347_185 ;
wire \top/processor/sha_core/n347_187 ;
wire \top/processor/sha_core/n347_189 ;
wire \top/processor/sha_core/n347_191 ;
wire \top/processor/sha_core/n347_193 ;
wire \top/processor/sha_core/n347_195 ;
wire \top/processor/sha_core/n348_165 ;
wire \top/processor/sha_core/n348_167 ;
wire \top/processor/sha_core/n348_169 ;
wire \top/processor/sha_core/n348_171 ;
wire \top/processor/sha_core/n348_173 ;
wire \top/processor/sha_core/n348_175 ;
wire \top/processor/sha_core/n348_177 ;
wire \top/processor/sha_core/n348_179 ;
wire \top/processor/sha_core/n348_181 ;
wire \top/processor/sha_core/n348_183 ;
wire \top/processor/sha_core/n348_185 ;
wire \top/processor/sha_core/n348_187 ;
wire \top/processor/sha_core/n348_189 ;
wire \top/processor/sha_core/n348_191 ;
wire \top/processor/sha_core/n348_193 ;
wire \top/processor/sha_core/n348_195 ;
wire \top/processor/sha_core/n349_165 ;
wire \top/processor/sha_core/n349_167 ;
wire \top/processor/sha_core/n349_169 ;
wire \top/processor/sha_core/n349_171 ;
wire \top/processor/sha_core/n349_173 ;
wire \top/processor/sha_core/n349_175 ;
wire \top/processor/sha_core/n349_177 ;
wire \top/processor/sha_core/n349_179 ;
wire \top/processor/sha_core/n349_181 ;
wire \top/processor/sha_core/n349_183 ;
wire \top/processor/sha_core/n349_185 ;
wire \top/processor/sha_core/n349_187 ;
wire \top/processor/sha_core/n349_189 ;
wire \top/processor/sha_core/n349_191 ;
wire \top/processor/sha_core/n349_193 ;
wire \top/processor/sha_core/n349_195 ;
wire \top/processor/sha_core/n350_165 ;
wire \top/processor/sha_core/n350_167 ;
wire \top/processor/sha_core/n350_169 ;
wire \top/processor/sha_core/n350_171 ;
wire \top/processor/sha_core/n350_173 ;
wire \top/processor/sha_core/n350_175 ;
wire \top/processor/sha_core/n350_177 ;
wire \top/processor/sha_core/n350_179 ;
wire \top/processor/sha_core/n350_181 ;
wire \top/processor/sha_core/n350_183 ;
wire \top/processor/sha_core/n350_185 ;
wire \top/processor/sha_core/n350_187 ;
wire \top/processor/sha_core/n350_189 ;
wire \top/processor/sha_core/n350_191 ;
wire \top/processor/sha_core/n350_193 ;
wire \top/processor/sha_core/n350_195 ;
wire \top/processor/sha_core/n351_165 ;
wire \top/processor/sha_core/n351_167 ;
wire \top/processor/sha_core/n351_169 ;
wire \top/processor/sha_core/n351_171 ;
wire \top/processor/sha_core/n351_173 ;
wire \top/processor/sha_core/n351_175 ;
wire \top/processor/sha_core/n351_177 ;
wire \top/processor/sha_core/n351_179 ;
wire \top/processor/sha_core/n351_181 ;
wire \top/processor/sha_core/n351_183 ;
wire \top/processor/sha_core/n351_185 ;
wire \top/processor/sha_core/n351_187 ;
wire \top/processor/sha_core/n351_189 ;
wire \top/processor/sha_core/n351_191 ;
wire \top/processor/sha_core/n351_193 ;
wire \top/processor/sha_core/n351_195 ;
wire \top/processor/sha_core/n352_165 ;
wire \top/processor/sha_core/n352_167 ;
wire \top/processor/sha_core/n352_169 ;
wire \top/processor/sha_core/n352_171 ;
wire \top/processor/sha_core/n352_173 ;
wire \top/processor/sha_core/n352_175 ;
wire \top/processor/sha_core/n352_177 ;
wire \top/processor/sha_core/n352_179 ;
wire \top/processor/sha_core/n352_181 ;
wire \top/processor/sha_core/n352_183 ;
wire \top/processor/sha_core/n352_185 ;
wire \top/processor/sha_core/n352_187 ;
wire \top/processor/sha_core/n352_189 ;
wire \top/processor/sha_core/n352_191 ;
wire \top/processor/sha_core/n352_193 ;
wire \top/processor/sha_core/n352_195 ;
wire \top/processor/sha_core/n353_165 ;
wire \top/processor/sha_core/n353_167 ;
wire \top/processor/sha_core/n353_169 ;
wire \top/processor/sha_core/n353_171 ;
wire \top/processor/sha_core/n353_173 ;
wire \top/processor/sha_core/n353_175 ;
wire \top/processor/sha_core/n353_177 ;
wire \top/processor/sha_core/n353_179 ;
wire \top/processor/sha_core/n353_181 ;
wire \top/processor/sha_core/n353_183 ;
wire \top/processor/sha_core/n353_185 ;
wire \top/processor/sha_core/n353_187 ;
wire \top/processor/sha_core/n353_189 ;
wire \top/processor/sha_core/n353_191 ;
wire \top/processor/sha_core/n353_193 ;
wire \top/processor/sha_core/n353_195 ;
wire \top/processor/sha_core/n354_165 ;
wire \top/processor/sha_core/n354_167 ;
wire \top/processor/sha_core/n354_169 ;
wire \top/processor/sha_core/n354_171 ;
wire \top/processor/sha_core/n354_173 ;
wire \top/processor/sha_core/n354_175 ;
wire \top/processor/sha_core/n354_177 ;
wire \top/processor/sha_core/n354_179 ;
wire \top/processor/sha_core/n354_181 ;
wire \top/processor/sha_core/n354_183 ;
wire \top/processor/sha_core/n354_185 ;
wire \top/processor/sha_core/n354_187 ;
wire \top/processor/sha_core/n354_189 ;
wire \top/processor/sha_core/n354_191 ;
wire \top/processor/sha_core/n354_193 ;
wire \top/processor/sha_core/n354_195 ;
wire \top/processor/sha_core/n355_165 ;
wire \top/processor/sha_core/n355_167 ;
wire \top/processor/sha_core/n355_169 ;
wire \top/processor/sha_core/n355_171 ;
wire \top/processor/sha_core/n355_173 ;
wire \top/processor/sha_core/n355_175 ;
wire \top/processor/sha_core/n355_177 ;
wire \top/processor/sha_core/n355_179 ;
wire \top/processor/sha_core/n355_181 ;
wire \top/processor/sha_core/n355_183 ;
wire \top/processor/sha_core/n355_185 ;
wire \top/processor/sha_core/n355_187 ;
wire \top/processor/sha_core/n355_189 ;
wire \top/processor/sha_core/n355_191 ;
wire \top/processor/sha_core/n355_193 ;
wire \top/processor/sha_core/n355_195 ;
wire \top/processor/sha_core/n356_165 ;
wire \top/processor/sha_core/n356_167 ;
wire \top/processor/sha_core/n356_169 ;
wire \top/processor/sha_core/n356_171 ;
wire \top/processor/sha_core/n356_173 ;
wire \top/processor/sha_core/n356_175 ;
wire \top/processor/sha_core/n356_177 ;
wire \top/processor/sha_core/n356_179 ;
wire \top/processor/sha_core/n356_181 ;
wire \top/processor/sha_core/n356_183 ;
wire \top/processor/sha_core/n356_185 ;
wire \top/processor/sha_core/n356_187 ;
wire \top/processor/sha_core/n356_189 ;
wire \top/processor/sha_core/n356_191 ;
wire \top/processor/sha_core/n356_193 ;
wire \top/processor/sha_core/n356_195 ;
wire \top/processor/sha_core/n357_165 ;
wire \top/processor/sha_core/n357_167 ;
wire \top/processor/sha_core/n357_169 ;
wire \top/processor/sha_core/n357_171 ;
wire \top/processor/sha_core/n357_173 ;
wire \top/processor/sha_core/n357_175 ;
wire \top/processor/sha_core/n357_177 ;
wire \top/processor/sha_core/n357_179 ;
wire \top/processor/sha_core/n357_181 ;
wire \top/processor/sha_core/n357_183 ;
wire \top/processor/sha_core/n357_185 ;
wire \top/processor/sha_core/n357_187 ;
wire \top/processor/sha_core/n357_189 ;
wire \top/processor/sha_core/n357_191 ;
wire \top/processor/sha_core/n357_193 ;
wire \top/processor/sha_core/n357_195 ;
wire \top/processor/sha_core/n358_165 ;
wire \top/processor/sha_core/n358_167 ;
wire \top/processor/sha_core/n358_169 ;
wire \top/processor/sha_core/n358_171 ;
wire \top/processor/sha_core/n358_173 ;
wire \top/processor/sha_core/n358_175 ;
wire \top/processor/sha_core/n358_177 ;
wire \top/processor/sha_core/n358_179 ;
wire \top/processor/sha_core/n358_181 ;
wire \top/processor/sha_core/n358_183 ;
wire \top/processor/sha_core/n358_185 ;
wire \top/processor/sha_core/n358_187 ;
wire \top/processor/sha_core/n358_189 ;
wire \top/processor/sha_core/n358_191 ;
wire \top/processor/sha_core/n358_193 ;
wire \top/processor/sha_core/n358_195 ;
wire \top/processor/sha_core/n3488_181 ;
wire \top/processor/sha_core/n3488_183 ;
wire \top/processor/sha_core/n3488_185 ;
wire \top/processor/sha_core/n3488_187 ;
wire \top/processor/sha_core/n3489_181 ;
wire \top/processor/sha_core/n3489_183 ;
wire \top/processor/sha_core/n3489_185 ;
wire \top/processor/sha_core/n3489_187 ;
wire \top/processor/sha_core/n3490_181 ;
wire \top/processor/sha_core/n3490_183 ;
wire \top/processor/sha_core/n3490_185 ;
wire \top/processor/sha_core/n3490_187 ;
wire \top/processor/sha_core/n3491_181 ;
wire \top/processor/sha_core/n3491_183 ;
wire \top/processor/sha_core/n3491_185 ;
wire \top/processor/sha_core/n3491_187 ;
wire \top/processor/sha_core/n3492_181 ;
wire \top/processor/sha_core/n3492_183 ;
wire \top/processor/sha_core/n3492_185 ;
wire \top/processor/sha_core/n3492_187 ;
wire \top/processor/sha_core/n3493_181 ;
wire \top/processor/sha_core/n3493_183 ;
wire \top/processor/sha_core/n3493_185 ;
wire \top/processor/sha_core/n3493_187 ;
wire \top/processor/sha_core/n3494_182 ;
wire \top/processor/sha_core/n3494_184 ;
wire \top/processor/sha_core/n3494_186 ;
wire \top/processor/sha_core/n3494_188 ;
wire \top/processor/sha_core/n3495_181 ;
wire \top/processor/sha_core/n3495_183 ;
wire \top/processor/sha_core/n3495_185 ;
wire \top/processor/sha_core/n3495_187 ;
wire \top/processor/sha_core/n3496_181 ;
wire \top/processor/sha_core/n3496_183 ;
wire \top/processor/sha_core/n3496_185 ;
wire \top/processor/sha_core/n3496_187 ;
wire \top/processor/sha_core/n3497_181 ;
wire \top/processor/sha_core/n3497_183 ;
wire \top/processor/sha_core/n3497_185 ;
wire \top/processor/sha_core/n3497_187 ;
wire \top/processor/sha_core/n3498_181 ;
wire \top/processor/sha_core/n3498_183 ;
wire \top/processor/sha_core/n3498_185 ;
wire \top/processor/sha_core/n3498_187 ;
wire \top/processor/sha_core/n3499_181 ;
wire \top/processor/sha_core/n3499_183 ;
wire \top/processor/sha_core/n3499_185 ;
wire \top/processor/sha_core/n3499_187 ;
wire \top/processor/sha_core/n3500_181 ;
wire \top/processor/sha_core/n3500_183 ;
wire \top/processor/sha_core/n3500_185 ;
wire \top/processor/sha_core/n3500_187 ;
wire \top/processor/sha_core/n3501_181 ;
wire \top/processor/sha_core/n3501_183 ;
wire \top/processor/sha_core/n3501_185 ;
wire \top/processor/sha_core/n3501_187 ;
wire \top/processor/sha_core/n3502_181 ;
wire \top/processor/sha_core/n3502_183 ;
wire \top/processor/sha_core/n3502_185 ;
wire \top/processor/sha_core/n3502_187 ;
wire \top/processor/sha_core/n3503_181 ;
wire \top/processor/sha_core/n3503_183 ;
wire \top/processor/sha_core/n3503_185 ;
wire \top/processor/sha_core/n3503_187 ;
wire \top/processor/sha_core/n3504_181 ;
wire \top/processor/sha_core/n3504_183 ;
wire \top/processor/sha_core/n3504_185 ;
wire \top/processor/sha_core/n3504_187 ;
wire \top/processor/sha_core/n3505_181 ;
wire \top/processor/sha_core/n3505_183 ;
wire \top/processor/sha_core/n3505_185 ;
wire \top/processor/sha_core/n3505_187 ;
wire \top/processor/sha_core/n3506_181 ;
wire \top/processor/sha_core/n3506_183 ;
wire \top/processor/sha_core/n3506_185 ;
wire \top/processor/sha_core/n3506_187 ;
wire \top/processor/sha_core/n3507_181 ;
wire \top/processor/sha_core/n3507_183 ;
wire \top/processor/sha_core/n3507_185 ;
wire \top/processor/sha_core/n3507_187 ;
wire \top/processor/sha_core/n3508_181 ;
wire \top/processor/sha_core/n3508_183 ;
wire \top/processor/sha_core/n3508_185 ;
wire \top/processor/sha_core/n3508_187 ;
wire \top/processor/sha_core/n3509_181 ;
wire \top/processor/sha_core/n3509_183 ;
wire \top/processor/sha_core/n3509_185 ;
wire \top/processor/sha_core/n3509_187 ;
wire \top/processor/sha_core/n3510_181 ;
wire \top/processor/sha_core/n3510_183 ;
wire \top/processor/sha_core/n3510_185 ;
wire \top/processor/sha_core/n3510_187 ;
wire \top/processor/sha_core/n3511_181 ;
wire \top/processor/sha_core/n3511_183 ;
wire \top/processor/sha_core/n3511_185 ;
wire \top/processor/sha_core/n3511_187 ;
wire \top/processor/sha_core/n3512_181 ;
wire \top/processor/sha_core/n3512_183 ;
wire \top/processor/sha_core/n3512_185 ;
wire \top/processor/sha_core/n3512_187 ;
wire \top/processor/sha_core/n3513_181 ;
wire \top/processor/sha_core/n3513_183 ;
wire \top/processor/sha_core/n3513_185 ;
wire \top/processor/sha_core/n3513_187 ;
wire \top/processor/sha_core/n3514_181 ;
wire \top/processor/sha_core/n3514_183 ;
wire \top/processor/sha_core/n3514_185 ;
wire \top/processor/sha_core/n3514_187 ;
wire \top/processor/sha_core/n3515_181 ;
wire \top/processor/sha_core/n3515_183 ;
wire \top/processor/sha_core/n3515_185 ;
wire \top/processor/sha_core/n3515_187 ;
wire \top/processor/sha_core/n3516_181 ;
wire \top/processor/sha_core/n3516_183 ;
wire \top/processor/sha_core/n3516_185 ;
wire \top/processor/sha_core/n3516_187 ;
wire \top/processor/sha_core/n3517_181 ;
wire \top/processor/sha_core/n3517_183 ;
wire \top/processor/sha_core/n3517_185 ;
wire \top/processor/sha_core/n3517_187 ;
wire \top/processor/sha_core/n3518_181 ;
wire \top/processor/sha_core/n3518_183 ;
wire \top/processor/sha_core/n3518_185 ;
wire \top/processor/sha_core/n3518_187 ;
wire \top/processor/sha_core/n3519_181 ;
wire \top/processor/sha_core/n3519_183 ;
wire \top/processor/sha_core/n3519_185 ;
wire \top/processor/sha_core/n3519_187 ;
wire \top/processor/sha_core/n3705_133 ;
wire \top/processor/sha_core/n3705_135 ;
wire \top/processor/sha_core/n3705_137 ;
wire \top/processor/sha_core/n3705_139 ;
wire \top/processor/sha_core/n3705_141 ;
wire \top/processor/sha_core/n3705_143 ;
wire \top/processor/sha_core/n3705_145 ;
wire \top/processor/sha_core/n3705_147 ;
wire \top/processor/sha_core/n3706_133 ;
wire \top/processor/sha_core/n3706_135 ;
wire \top/processor/sha_core/n3706_137 ;
wire \top/processor/sha_core/n3706_139 ;
wire \top/processor/sha_core/n3706_141 ;
wire \top/processor/sha_core/n3706_143 ;
wire \top/processor/sha_core/n3706_145 ;
wire \top/processor/sha_core/n3706_147 ;
wire \top/processor/sha_core/n3707_133 ;
wire \top/processor/sha_core/n3707_135 ;
wire \top/processor/sha_core/n3707_137 ;
wire \top/processor/sha_core/n3707_139 ;
wire \top/processor/sha_core/n3707_141 ;
wire \top/processor/sha_core/n3707_143 ;
wire \top/processor/sha_core/n3707_145 ;
wire \top/processor/sha_core/n3707_147 ;
wire \top/processor/sha_core/n3708_133 ;
wire \top/processor/sha_core/n3708_135 ;
wire \top/processor/sha_core/n3708_137 ;
wire \top/processor/sha_core/n3708_139 ;
wire \top/processor/sha_core/n3708_141 ;
wire \top/processor/sha_core/n3708_143 ;
wire \top/processor/sha_core/n3708_145 ;
wire \top/processor/sha_core/n3708_147 ;
wire \top/processor/sha_core/n3709_133 ;
wire \top/processor/sha_core/n3709_135 ;
wire \top/processor/sha_core/n3709_137 ;
wire \top/processor/sha_core/n3709_139 ;
wire \top/processor/sha_core/n3709_141 ;
wire \top/processor/sha_core/n3709_143 ;
wire \top/processor/sha_core/n3709_145 ;
wire \top/processor/sha_core/n3709_147 ;
wire \top/processor/sha_core/n3710_133 ;
wire \top/processor/sha_core/n3710_135 ;
wire \top/processor/sha_core/n3710_137 ;
wire \top/processor/sha_core/n3710_139 ;
wire \top/processor/sha_core/n3710_141 ;
wire \top/processor/sha_core/n3710_143 ;
wire \top/processor/sha_core/n3710_145 ;
wire \top/processor/sha_core/n3710_147 ;
wire \top/processor/sha_core/n3711_133 ;
wire \top/processor/sha_core/n3711_135 ;
wire \top/processor/sha_core/n3711_137 ;
wire \top/processor/sha_core/n3711_139 ;
wire \top/processor/sha_core/n3711_141 ;
wire \top/processor/sha_core/n3711_143 ;
wire \top/processor/sha_core/n3711_145 ;
wire \top/processor/sha_core/n3711_147 ;
wire \top/processor/sha_core/n3712_133 ;
wire \top/processor/sha_core/n3712_135 ;
wire \top/processor/sha_core/n3712_137 ;
wire \top/processor/sha_core/n3712_139 ;
wire \top/processor/sha_core/n3712_141 ;
wire \top/processor/sha_core/n3712_143 ;
wire \top/processor/sha_core/n3712_145 ;
wire \top/processor/sha_core/n3712_147 ;
wire \top/processor/sha_core/n3713_133 ;
wire \top/processor/sha_core/n3713_135 ;
wire \top/processor/sha_core/n3713_137 ;
wire \top/processor/sha_core/n3713_139 ;
wire \top/processor/sha_core/n3713_141 ;
wire \top/processor/sha_core/n3713_143 ;
wire \top/processor/sha_core/n3713_145 ;
wire \top/processor/sha_core/n3713_147 ;
wire \top/processor/sha_core/n3714_133 ;
wire \top/processor/sha_core/n3714_135 ;
wire \top/processor/sha_core/n3714_137 ;
wire \top/processor/sha_core/n3714_139 ;
wire \top/processor/sha_core/n3714_141 ;
wire \top/processor/sha_core/n3714_143 ;
wire \top/processor/sha_core/n3714_145 ;
wire \top/processor/sha_core/n3714_147 ;
wire \top/processor/sha_core/n3715_133 ;
wire \top/processor/sha_core/n3715_135 ;
wire \top/processor/sha_core/n3715_137 ;
wire \top/processor/sha_core/n3715_139 ;
wire \top/processor/sha_core/n3715_141 ;
wire \top/processor/sha_core/n3715_143 ;
wire \top/processor/sha_core/n3715_145 ;
wire \top/processor/sha_core/n3715_147 ;
wire \top/processor/sha_core/n3716_133 ;
wire \top/processor/sha_core/n3716_135 ;
wire \top/processor/sha_core/n3716_137 ;
wire \top/processor/sha_core/n3716_139 ;
wire \top/processor/sha_core/n3716_141 ;
wire \top/processor/sha_core/n3716_143 ;
wire \top/processor/sha_core/n3716_145 ;
wire \top/processor/sha_core/n3716_147 ;
wire \top/processor/sha_core/n3717_133 ;
wire \top/processor/sha_core/n3717_135 ;
wire \top/processor/sha_core/n3717_137 ;
wire \top/processor/sha_core/n3717_139 ;
wire \top/processor/sha_core/n3717_141 ;
wire \top/processor/sha_core/n3717_143 ;
wire \top/processor/sha_core/n3717_145 ;
wire \top/processor/sha_core/n3717_147 ;
wire \top/processor/sha_core/n3718_133 ;
wire \top/processor/sha_core/n3718_135 ;
wire \top/processor/sha_core/n3718_137 ;
wire \top/processor/sha_core/n3718_139 ;
wire \top/processor/sha_core/n3718_141 ;
wire \top/processor/sha_core/n3718_143 ;
wire \top/processor/sha_core/n3718_145 ;
wire \top/processor/sha_core/n3718_147 ;
wire \top/processor/sha_core/n3719_133 ;
wire \top/processor/sha_core/n3719_135 ;
wire \top/processor/sha_core/n3719_137 ;
wire \top/processor/sha_core/n3719_139 ;
wire \top/processor/sha_core/n3719_141 ;
wire \top/processor/sha_core/n3719_143 ;
wire \top/processor/sha_core/n3719_145 ;
wire \top/processor/sha_core/n3719_147 ;
wire \top/processor/sha_core/n3720_133 ;
wire \top/processor/sha_core/n3720_135 ;
wire \top/processor/sha_core/n3720_137 ;
wire \top/processor/sha_core/n3720_139 ;
wire \top/processor/sha_core/n3720_141 ;
wire \top/processor/sha_core/n3720_143 ;
wire \top/processor/sha_core/n3720_145 ;
wire \top/processor/sha_core/n3720_147 ;
wire \top/processor/sha_core/n3721_133 ;
wire \top/processor/sha_core/n3721_135 ;
wire \top/processor/sha_core/n3721_137 ;
wire \top/processor/sha_core/n3721_139 ;
wire \top/processor/sha_core/n3721_141 ;
wire \top/processor/sha_core/n3721_143 ;
wire \top/processor/sha_core/n3721_145 ;
wire \top/processor/sha_core/n3721_147 ;
wire \top/processor/sha_core/n3722_133 ;
wire \top/processor/sha_core/n3722_135 ;
wire \top/processor/sha_core/n3722_137 ;
wire \top/processor/sha_core/n3722_139 ;
wire \top/processor/sha_core/n3722_141 ;
wire \top/processor/sha_core/n3722_143 ;
wire \top/processor/sha_core/n3722_145 ;
wire \top/processor/sha_core/n3722_147 ;
wire \top/processor/sha_core/n3723_133 ;
wire \top/processor/sha_core/n3723_135 ;
wire \top/processor/sha_core/n3723_137 ;
wire \top/processor/sha_core/n3723_139 ;
wire \top/processor/sha_core/n3723_141 ;
wire \top/processor/sha_core/n3723_143 ;
wire \top/processor/sha_core/n3723_145 ;
wire \top/processor/sha_core/n3723_147 ;
wire \top/processor/sha_core/n3724_133 ;
wire \top/processor/sha_core/n3724_135 ;
wire \top/processor/sha_core/n3724_137 ;
wire \top/processor/sha_core/n3724_139 ;
wire \top/processor/sha_core/n3724_141 ;
wire \top/processor/sha_core/n3724_143 ;
wire \top/processor/sha_core/n3724_145 ;
wire \top/processor/sha_core/n3724_147 ;
wire \top/processor/sha_core/n3725_133 ;
wire \top/processor/sha_core/n3725_135 ;
wire \top/processor/sha_core/n3725_137 ;
wire \top/processor/sha_core/n3725_139 ;
wire \top/processor/sha_core/n3725_141 ;
wire \top/processor/sha_core/n3725_143 ;
wire \top/processor/sha_core/n3725_145 ;
wire \top/processor/sha_core/n3725_147 ;
wire \top/processor/sha_core/n3726_133 ;
wire \top/processor/sha_core/n3726_135 ;
wire \top/processor/sha_core/n3726_137 ;
wire \top/processor/sha_core/n3726_139 ;
wire \top/processor/sha_core/n3726_141 ;
wire \top/processor/sha_core/n3726_143 ;
wire \top/processor/sha_core/n3726_145 ;
wire \top/processor/sha_core/n3726_147 ;
wire \top/processor/sha_core/n3727_133 ;
wire \top/processor/sha_core/n3727_135 ;
wire \top/processor/sha_core/n3727_137 ;
wire \top/processor/sha_core/n3727_139 ;
wire \top/processor/sha_core/n3727_141 ;
wire \top/processor/sha_core/n3727_143 ;
wire \top/processor/sha_core/n3727_145 ;
wire \top/processor/sha_core/n3727_147 ;
wire \top/processor/sha_core/n3728_133 ;
wire \top/processor/sha_core/n3728_135 ;
wire \top/processor/sha_core/n3728_137 ;
wire \top/processor/sha_core/n3728_139 ;
wire \top/processor/sha_core/n3728_141 ;
wire \top/processor/sha_core/n3728_143 ;
wire \top/processor/sha_core/n3728_145 ;
wire \top/processor/sha_core/n3728_147 ;
wire \top/processor/sha_core/n3729_133 ;
wire \top/processor/sha_core/n3729_135 ;
wire \top/processor/sha_core/n3729_137 ;
wire \top/processor/sha_core/n3729_139 ;
wire \top/processor/sha_core/n3729_141 ;
wire \top/processor/sha_core/n3729_143 ;
wire \top/processor/sha_core/n3729_145 ;
wire \top/processor/sha_core/n3729_147 ;
wire \top/processor/sha_core/n3730_133 ;
wire \top/processor/sha_core/n3730_135 ;
wire \top/processor/sha_core/n3730_137 ;
wire \top/processor/sha_core/n3730_139 ;
wire \top/processor/sha_core/n3730_141 ;
wire \top/processor/sha_core/n3730_143 ;
wire \top/processor/sha_core/n3730_145 ;
wire \top/processor/sha_core/n3730_147 ;
wire \top/processor/sha_core/n3731_133 ;
wire \top/processor/sha_core/n3731_135 ;
wire \top/processor/sha_core/n3731_137 ;
wire \top/processor/sha_core/n3731_139 ;
wire \top/processor/sha_core/n3731_141 ;
wire \top/processor/sha_core/n3731_143 ;
wire \top/processor/sha_core/n3731_145 ;
wire \top/processor/sha_core/n3731_147 ;
wire \top/processor/sha_core/n3732_133 ;
wire \top/processor/sha_core/n3732_135 ;
wire \top/processor/sha_core/n3732_137 ;
wire \top/processor/sha_core/n3732_139 ;
wire \top/processor/sha_core/n3732_141 ;
wire \top/processor/sha_core/n3732_143 ;
wire \top/processor/sha_core/n3732_145 ;
wire \top/processor/sha_core/n3732_147 ;
wire \top/processor/sha_core/n3733_133 ;
wire \top/processor/sha_core/n3733_135 ;
wire \top/processor/sha_core/n3733_137 ;
wire \top/processor/sha_core/n3733_139 ;
wire \top/processor/sha_core/n3733_141 ;
wire \top/processor/sha_core/n3733_143 ;
wire \top/processor/sha_core/n3733_145 ;
wire \top/processor/sha_core/n3733_147 ;
wire \top/processor/sha_core/n3734_133 ;
wire \top/processor/sha_core/n3734_135 ;
wire \top/processor/sha_core/n3734_137 ;
wire \top/processor/sha_core/n3734_139 ;
wire \top/processor/sha_core/n3734_141 ;
wire \top/processor/sha_core/n3734_143 ;
wire \top/processor/sha_core/n3734_145 ;
wire \top/processor/sha_core/n3734_147 ;
wire \top/processor/sha_core/n3735_133 ;
wire \top/processor/sha_core/n3735_135 ;
wire \top/processor/sha_core/n3735_137 ;
wire \top/processor/sha_core/n3735_139 ;
wire \top/processor/sha_core/n3735_141 ;
wire \top/processor/sha_core/n3735_143 ;
wire \top/processor/sha_core/n3735_145 ;
wire \top/processor/sha_core/n3735_147 ;
wire \top/processor/sha_core/n3736_133 ;
wire \top/processor/sha_core/n3736_135 ;
wire \top/processor/sha_core/n3736_137 ;
wire \top/processor/sha_core/n3736_139 ;
wire \top/processor/sha_core/n3736_141 ;
wire \top/processor/sha_core/n3736_143 ;
wire \top/processor/sha_core/n3736_145 ;
wire \top/processor/sha_core/n3736_147 ;
wire \top/processor/sha_core/n3860_133 ;
wire \top/processor/sha_core/n3860_135 ;
wire \top/processor/sha_core/n3860_137 ;
wire \top/processor/sha_core/n3860_139 ;
wire \top/processor/sha_core/n3861_133 ;
wire \top/processor/sha_core/n3861_135 ;
wire \top/processor/sha_core/n3861_137 ;
wire \top/processor/sha_core/n3861_139 ;
wire \top/processor/sha_core/n3862_133 ;
wire \top/processor/sha_core/n3862_135 ;
wire \top/processor/sha_core/n3862_137 ;
wire \top/processor/sha_core/n3862_139 ;
wire \top/processor/sha_core/n3863_133 ;
wire \top/processor/sha_core/n3863_135 ;
wire \top/processor/sha_core/n3863_137 ;
wire \top/processor/sha_core/n3863_139 ;
wire \top/processor/sha_core/n3864_133 ;
wire \top/processor/sha_core/n3864_135 ;
wire \top/processor/sha_core/n3864_137 ;
wire \top/processor/sha_core/n3864_139 ;
wire \top/processor/sha_core/n3865_133 ;
wire \top/processor/sha_core/n3865_135 ;
wire \top/processor/sha_core/n3865_137 ;
wire \top/processor/sha_core/n3865_139 ;
wire \top/processor/sha_core/n3866_133 ;
wire \top/processor/sha_core/n3866_135 ;
wire \top/processor/sha_core/n3866_137 ;
wire \top/processor/sha_core/n3866_139 ;
wire \top/processor/sha_core/n3867_133 ;
wire \top/processor/sha_core/n3867_135 ;
wire \top/processor/sha_core/n3867_137 ;
wire \top/processor/sha_core/n3867_139 ;
wire \top/processor/sha_core/n3868_133 ;
wire \top/processor/sha_core/n3868_135 ;
wire \top/processor/sha_core/n3868_137 ;
wire \top/processor/sha_core/n3868_139 ;
wire \top/processor/sha_core/n3869_133 ;
wire \top/processor/sha_core/n3869_135 ;
wire \top/processor/sha_core/n3869_137 ;
wire \top/processor/sha_core/n3869_139 ;
wire \top/processor/sha_core/n3870_133 ;
wire \top/processor/sha_core/n3870_135 ;
wire \top/processor/sha_core/n3870_137 ;
wire \top/processor/sha_core/n3870_139 ;
wire \top/processor/sha_core/n3871_133 ;
wire \top/processor/sha_core/n3871_135 ;
wire \top/processor/sha_core/n3871_137 ;
wire \top/processor/sha_core/n3871_139 ;
wire \top/processor/sha_core/n3872_133 ;
wire \top/processor/sha_core/n3872_135 ;
wire \top/processor/sha_core/n3872_137 ;
wire \top/processor/sha_core/n3872_139 ;
wire \top/processor/sha_core/n3873_133 ;
wire \top/processor/sha_core/n3873_135 ;
wire \top/processor/sha_core/n3873_137 ;
wire \top/processor/sha_core/n3873_139 ;
wire \top/processor/sha_core/n3874_133 ;
wire \top/processor/sha_core/n3874_135 ;
wire \top/processor/sha_core/n3874_137 ;
wire \top/processor/sha_core/n3874_139 ;
wire \top/processor/sha_core/n3875_133 ;
wire \top/processor/sha_core/n3875_135 ;
wire \top/processor/sha_core/n3875_137 ;
wire \top/processor/sha_core/n3875_139 ;
wire \top/processor/sha_core/n3876_133 ;
wire \top/processor/sha_core/n3876_135 ;
wire \top/processor/sha_core/n3876_137 ;
wire \top/processor/sha_core/n3876_139 ;
wire \top/processor/sha_core/n3877_133 ;
wire \top/processor/sha_core/n3877_135 ;
wire \top/processor/sha_core/n3877_137 ;
wire \top/processor/sha_core/n3877_139 ;
wire \top/processor/sha_core/n3878_133 ;
wire \top/processor/sha_core/n3878_135 ;
wire \top/processor/sha_core/n3878_137 ;
wire \top/processor/sha_core/n3878_139 ;
wire \top/processor/sha_core/n3879_133 ;
wire \top/processor/sha_core/n3879_135 ;
wire \top/processor/sha_core/n3879_137 ;
wire \top/processor/sha_core/n3879_139 ;
wire \top/processor/sha_core/n3880_133 ;
wire \top/processor/sha_core/n3880_135 ;
wire \top/processor/sha_core/n3880_137 ;
wire \top/processor/sha_core/n3880_139 ;
wire \top/processor/sha_core/n3881_133 ;
wire \top/processor/sha_core/n3881_135 ;
wire \top/processor/sha_core/n3881_137 ;
wire \top/processor/sha_core/n3881_139 ;
wire \top/processor/sha_core/n3882_133 ;
wire \top/processor/sha_core/n3882_135 ;
wire \top/processor/sha_core/n3882_137 ;
wire \top/processor/sha_core/n3882_139 ;
wire \top/processor/sha_core/n3883_133 ;
wire \top/processor/sha_core/n3883_135 ;
wire \top/processor/sha_core/n3883_137 ;
wire \top/processor/sha_core/n3883_139 ;
wire \top/processor/sha_core/n3884_133 ;
wire \top/processor/sha_core/n3884_135 ;
wire \top/processor/sha_core/n3884_137 ;
wire \top/processor/sha_core/n3884_139 ;
wire \top/processor/sha_core/n3885_133 ;
wire \top/processor/sha_core/n3885_135 ;
wire \top/processor/sha_core/n3885_137 ;
wire \top/processor/sha_core/n3885_139 ;
wire \top/processor/sha_core/n3886_133 ;
wire \top/processor/sha_core/n3886_135 ;
wire \top/processor/sha_core/n3886_137 ;
wire \top/processor/sha_core/n3886_139 ;
wire \top/processor/sha_core/n3887_133 ;
wire \top/processor/sha_core/n3887_135 ;
wire \top/processor/sha_core/n3887_137 ;
wire \top/processor/sha_core/n3887_139 ;
wire \top/processor/sha_core/n3888_133 ;
wire \top/processor/sha_core/n3888_135 ;
wire \top/processor/sha_core/n3888_137 ;
wire \top/processor/sha_core/n3888_139 ;
wire \top/processor/sha_core/n3889_133 ;
wire \top/processor/sha_core/n3889_135 ;
wire \top/processor/sha_core/n3889_137 ;
wire \top/processor/sha_core/n3889_139 ;
wire \top/processor/sha_core/n3890_133 ;
wire \top/processor/sha_core/n3890_135 ;
wire \top/processor/sha_core/n3890_137 ;
wire \top/processor/sha_core/n3890_139 ;
wire \top/processor/sha_core/n3891_133 ;
wire \top/processor/sha_core/n3891_135 ;
wire \top/processor/sha_core/n3891_137 ;
wire \top/processor/sha_core/n3891_139 ;
wire \top/processor/sha_core/n327_197 ;
wire \top/processor/sha_core/n327_199 ;
wire \top/processor/sha_core/n327_201 ;
wire \top/processor/sha_core/n327_203 ;
wire \top/processor/sha_core/n327_205 ;
wire \top/processor/sha_core/n327_207 ;
wire \top/processor/sha_core/n327_209 ;
wire \top/processor/sha_core/n327_211 ;
wire \top/processor/sha_core/n328_197 ;
wire \top/processor/sha_core/n328_199 ;
wire \top/processor/sha_core/n328_201 ;
wire \top/processor/sha_core/n328_203 ;
wire \top/processor/sha_core/n328_205 ;
wire \top/processor/sha_core/n328_207 ;
wire \top/processor/sha_core/n328_209 ;
wire \top/processor/sha_core/n328_211 ;
wire \top/processor/sha_core/n329_197 ;
wire \top/processor/sha_core/n329_199 ;
wire \top/processor/sha_core/n329_201 ;
wire \top/processor/sha_core/n329_203 ;
wire \top/processor/sha_core/n329_205 ;
wire \top/processor/sha_core/n329_207 ;
wire \top/processor/sha_core/n329_209 ;
wire \top/processor/sha_core/n329_211 ;
wire \top/processor/sha_core/n330_197 ;
wire \top/processor/sha_core/n330_199 ;
wire \top/processor/sha_core/n330_201 ;
wire \top/processor/sha_core/n330_203 ;
wire \top/processor/sha_core/n330_205 ;
wire \top/processor/sha_core/n330_207 ;
wire \top/processor/sha_core/n330_209 ;
wire \top/processor/sha_core/n330_211 ;
wire \top/processor/sha_core/n331_197 ;
wire \top/processor/sha_core/n331_199 ;
wire \top/processor/sha_core/n331_201 ;
wire \top/processor/sha_core/n331_203 ;
wire \top/processor/sha_core/n331_205 ;
wire \top/processor/sha_core/n331_207 ;
wire \top/processor/sha_core/n331_209 ;
wire \top/processor/sha_core/n331_211 ;
wire \top/processor/sha_core/n332_197 ;
wire \top/processor/sha_core/n332_199 ;
wire \top/processor/sha_core/n332_201 ;
wire \top/processor/sha_core/n332_203 ;
wire \top/processor/sha_core/n332_205 ;
wire \top/processor/sha_core/n332_207 ;
wire \top/processor/sha_core/n332_209 ;
wire \top/processor/sha_core/n332_211 ;
wire \top/processor/sha_core/n333_197 ;
wire \top/processor/sha_core/n333_199 ;
wire \top/processor/sha_core/n333_201 ;
wire \top/processor/sha_core/n333_203 ;
wire \top/processor/sha_core/n333_205 ;
wire \top/processor/sha_core/n333_207 ;
wire \top/processor/sha_core/n333_209 ;
wire \top/processor/sha_core/n333_211 ;
wire \top/processor/sha_core/n334_197 ;
wire \top/processor/sha_core/n334_199 ;
wire \top/processor/sha_core/n334_201 ;
wire \top/processor/sha_core/n334_203 ;
wire \top/processor/sha_core/n334_205 ;
wire \top/processor/sha_core/n334_207 ;
wire \top/processor/sha_core/n334_209 ;
wire \top/processor/sha_core/n334_211 ;
wire \top/processor/sha_core/n335_197 ;
wire \top/processor/sha_core/n335_199 ;
wire \top/processor/sha_core/n335_201 ;
wire \top/processor/sha_core/n335_203 ;
wire \top/processor/sha_core/n335_205 ;
wire \top/processor/sha_core/n335_207 ;
wire \top/processor/sha_core/n335_209 ;
wire \top/processor/sha_core/n335_211 ;
wire \top/processor/sha_core/n336_197 ;
wire \top/processor/sha_core/n336_199 ;
wire \top/processor/sha_core/n336_201 ;
wire \top/processor/sha_core/n336_203 ;
wire \top/processor/sha_core/n336_205 ;
wire \top/processor/sha_core/n336_207 ;
wire \top/processor/sha_core/n336_209 ;
wire \top/processor/sha_core/n336_211 ;
wire \top/processor/sha_core/n337_197 ;
wire \top/processor/sha_core/n337_199 ;
wire \top/processor/sha_core/n337_201 ;
wire \top/processor/sha_core/n337_203 ;
wire \top/processor/sha_core/n337_205 ;
wire \top/processor/sha_core/n337_207 ;
wire \top/processor/sha_core/n337_209 ;
wire \top/processor/sha_core/n337_211 ;
wire \top/processor/sha_core/n338_197 ;
wire \top/processor/sha_core/n338_199 ;
wire \top/processor/sha_core/n338_201 ;
wire \top/processor/sha_core/n338_203 ;
wire \top/processor/sha_core/n338_205 ;
wire \top/processor/sha_core/n338_207 ;
wire \top/processor/sha_core/n338_209 ;
wire \top/processor/sha_core/n338_211 ;
wire \top/processor/sha_core/n339_197 ;
wire \top/processor/sha_core/n339_199 ;
wire \top/processor/sha_core/n339_201 ;
wire \top/processor/sha_core/n339_203 ;
wire \top/processor/sha_core/n339_205 ;
wire \top/processor/sha_core/n339_207 ;
wire \top/processor/sha_core/n339_209 ;
wire \top/processor/sha_core/n339_211 ;
wire \top/processor/sha_core/n340_197 ;
wire \top/processor/sha_core/n340_199 ;
wire \top/processor/sha_core/n340_201 ;
wire \top/processor/sha_core/n340_203 ;
wire \top/processor/sha_core/n340_205 ;
wire \top/processor/sha_core/n340_207 ;
wire \top/processor/sha_core/n340_209 ;
wire \top/processor/sha_core/n340_211 ;
wire \top/processor/sha_core/n341_197 ;
wire \top/processor/sha_core/n341_199 ;
wire \top/processor/sha_core/n341_201 ;
wire \top/processor/sha_core/n341_203 ;
wire \top/processor/sha_core/n341_205 ;
wire \top/processor/sha_core/n341_207 ;
wire \top/processor/sha_core/n341_209 ;
wire \top/processor/sha_core/n341_211 ;
wire \top/processor/sha_core/n342_197 ;
wire \top/processor/sha_core/n342_199 ;
wire \top/processor/sha_core/n342_201 ;
wire \top/processor/sha_core/n342_203 ;
wire \top/processor/sha_core/n342_205 ;
wire \top/processor/sha_core/n342_207 ;
wire \top/processor/sha_core/n342_209 ;
wire \top/processor/sha_core/n342_211 ;
wire \top/processor/sha_core/n343_197 ;
wire \top/processor/sha_core/n343_199 ;
wire \top/processor/sha_core/n343_201 ;
wire \top/processor/sha_core/n343_203 ;
wire \top/processor/sha_core/n343_205 ;
wire \top/processor/sha_core/n343_207 ;
wire \top/processor/sha_core/n343_209 ;
wire \top/processor/sha_core/n343_211 ;
wire \top/processor/sha_core/n344_197 ;
wire \top/processor/sha_core/n344_199 ;
wire \top/processor/sha_core/n344_201 ;
wire \top/processor/sha_core/n344_203 ;
wire \top/processor/sha_core/n344_205 ;
wire \top/processor/sha_core/n344_207 ;
wire \top/processor/sha_core/n344_209 ;
wire \top/processor/sha_core/n344_211 ;
wire \top/processor/sha_core/n345_197 ;
wire \top/processor/sha_core/n345_199 ;
wire \top/processor/sha_core/n345_201 ;
wire \top/processor/sha_core/n345_203 ;
wire \top/processor/sha_core/n345_205 ;
wire \top/processor/sha_core/n345_207 ;
wire \top/processor/sha_core/n345_209 ;
wire \top/processor/sha_core/n345_211 ;
wire \top/processor/sha_core/n346_197 ;
wire \top/processor/sha_core/n346_199 ;
wire \top/processor/sha_core/n346_201 ;
wire \top/processor/sha_core/n346_203 ;
wire \top/processor/sha_core/n346_205 ;
wire \top/processor/sha_core/n346_207 ;
wire \top/processor/sha_core/n346_209 ;
wire \top/processor/sha_core/n346_211 ;
wire \top/processor/sha_core/n347_197 ;
wire \top/processor/sha_core/n347_199 ;
wire \top/processor/sha_core/n347_201 ;
wire \top/processor/sha_core/n347_203 ;
wire \top/processor/sha_core/n347_205 ;
wire \top/processor/sha_core/n347_207 ;
wire \top/processor/sha_core/n347_209 ;
wire \top/processor/sha_core/n347_211 ;
wire \top/processor/sha_core/n348_197 ;
wire \top/processor/sha_core/n348_199 ;
wire \top/processor/sha_core/n348_201 ;
wire \top/processor/sha_core/n348_203 ;
wire \top/processor/sha_core/n348_205 ;
wire \top/processor/sha_core/n348_207 ;
wire \top/processor/sha_core/n348_209 ;
wire \top/processor/sha_core/n348_211 ;
wire \top/processor/sha_core/n349_197 ;
wire \top/processor/sha_core/n349_199 ;
wire \top/processor/sha_core/n349_201 ;
wire \top/processor/sha_core/n349_203 ;
wire \top/processor/sha_core/n349_205 ;
wire \top/processor/sha_core/n349_207 ;
wire \top/processor/sha_core/n349_209 ;
wire \top/processor/sha_core/n349_211 ;
wire \top/processor/sha_core/n350_197 ;
wire \top/processor/sha_core/n350_199 ;
wire \top/processor/sha_core/n350_201 ;
wire \top/processor/sha_core/n350_203 ;
wire \top/processor/sha_core/n350_205 ;
wire \top/processor/sha_core/n350_207 ;
wire \top/processor/sha_core/n350_209 ;
wire \top/processor/sha_core/n350_211 ;
wire \top/processor/sha_core/n351_197 ;
wire \top/processor/sha_core/n351_199 ;
wire \top/processor/sha_core/n351_201 ;
wire \top/processor/sha_core/n351_203 ;
wire \top/processor/sha_core/n351_205 ;
wire \top/processor/sha_core/n351_207 ;
wire \top/processor/sha_core/n351_209 ;
wire \top/processor/sha_core/n351_211 ;
wire \top/processor/sha_core/n352_197 ;
wire \top/processor/sha_core/n352_199 ;
wire \top/processor/sha_core/n352_201 ;
wire \top/processor/sha_core/n352_203 ;
wire \top/processor/sha_core/n352_205 ;
wire \top/processor/sha_core/n352_207 ;
wire \top/processor/sha_core/n352_209 ;
wire \top/processor/sha_core/n352_211 ;
wire \top/processor/sha_core/n353_197 ;
wire \top/processor/sha_core/n353_199 ;
wire \top/processor/sha_core/n353_201 ;
wire \top/processor/sha_core/n353_203 ;
wire \top/processor/sha_core/n353_205 ;
wire \top/processor/sha_core/n353_207 ;
wire \top/processor/sha_core/n353_209 ;
wire \top/processor/sha_core/n353_211 ;
wire \top/processor/sha_core/n354_197 ;
wire \top/processor/sha_core/n354_199 ;
wire \top/processor/sha_core/n354_201 ;
wire \top/processor/sha_core/n354_203 ;
wire \top/processor/sha_core/n354_205 ;
wire \top/processor/sha_core/n354_207 ;
wire \top/processor/sha_core/n354_209 ;
wire \top/processor/sha_core/n354_211 ;
wire \top/processor/sha_core/n355_197 ;
wire \top/processor/sha_core/n355_199 ;
wire \top/processor/sha_core/n355_201 ;
wire \top/processor/sha_core/n355_203 ;
wire \top/processor/sha_core/n355_205 ;
wire \top/processor/sha_core/n355_207 ;
wire \top/processor/sha_core/n355_209 ;
wire \top/processor/sha_core/n355_211 ;
wire \top/processor/sha_core/n356_197 ;
wire \top/processor/sha_core/n356_199 ;
wire \top/processor/sha_core/n356_201 ;
wire \top/processor/sha_core/n356_203 ;
wire \top/processor/sha_core/n356_205 ;
wire \top/processor/sha_core/n356_207 ;
wire \top/processor/sha_core/n356_209 ;
wire \top/processor/sha_core/n356_211 ;
wire \top/processor/sha_core/n357_197 ;
wire \top/processor/sha_core/n357_199 ;
wire \top/processor/sha_core/n357_201 ;
wire \top/processor/sha_core/n357_203 ;
wire \top/processor/sha_core/n357_205 ;
wire \top/processor/sha_core/n357_207 ;
wire \top/processor/sha_core/n357_209 ;
wire \top/processor/sha_core/n357_211 ;
wire \top/processor/sha_core/n358_197 ;
wire \top/processor/sha_core/n358_199 ;
wire \top/processor/sha_core/n358_201 ;
wire \top/processor/sha_core/n358_203 ;
wire \top/processor/sha_core/n358_205 ;
wire \top/processor/sha_core/n358_207 ;
wire \top/processor/sha_core/n358_209 ;
wire \top/processor/sha_core/n358_211 ;
wire \top/processor/sha_core/n3488_189 ;
wire \top/processor/sha_core/n3488_191 ;
wire \top/processor/sha_core/n3489_189 ;
wire \top/processor/sha_core/n3489_191 ;
wire \top/processor/sha_core/n3490_189 ;
wire \top/processor/sha_core/n3490_191 ;
wire \top/processor/sha_core/n3491_189 ;
wire \top/processor/sha_core/n3491_191 ;
wire \top/processor/sha_core/n3492_189 ;
wire \top/processor/sha_core/n3492_191 ;
wire \top/processor/sha_core/n3493_189 ;
wire \top/processor/sha_core/n3493_191 ;
wire \top/processor/sha_core/n3494_190 ;
wire \top/processor/sha_core/n3494_192 ;
wire \top/processor/sha_core/n3495_189 ;
wire \top/processor/sha_core/n3495_191 ;
wire \top/processor/sha_core/n3496_189 ;
wire \top/processor/sha_core/n3496_191 ;
wire \top/processor/sha_core/n3497_189 ;
wire \top/processor/sha_core/n3497_191 ;
wire \top/processor/sha_core/n3498_189 ;
wire \top/processor/sha_core/n3498_191 ;
wire \top/processor/sha_core/n3499_189 ;
wire \top/processor/sha_core/n3499_191 ;
wire \top/processor/sha_core/n3500_189 ;
wire \top/processor/sha_core/n3500_191 ;
wire \top/processor/sha_core/n3501_189 ;
wire \top/processor/sha_core/n3501_191 ;
wire \top/processor/sha_core/n3502_189 ;
wire \top/processor/sha_core/n3502_191 ;
wire \top/processor/sha_core/n3503_189 ;
wire \top/processor/sha_core/n3503_191 ;
wire \top/processor/sha_core/n3504_189 ;
wire \top/processor/sha_core/n3504_191 ;
wire \top/processor/sha_core/n3505_189 ;
wire \top/processor/sha_core/n3505_191 ;
wire \top/processor/sha_core/n3506_189 ;
wire \top/processor/sha_core/n3506_191 ;
wire \top/processor/sha_core/n3507_189 ;
wire \top/processor/sha_core/n3507_191 ;
wire \top/processor/sha_core/n3508_189 ;
wire \top/processor/sha_core/n3508_191 ;
wire \top/processor/sha_core/n3509_189 ;
wire \top/processor/sha_core/n3509_191 ;
wire \top/processor/sha_core/n3510_189 ;
wire \top/processor/sha_core/n3510_191 ;
wire \top/processor/sha_core/n3511_189 ;
wire \top/processor/sha_core/n3511_191 ;
wire \top/processor/sha_core/n3512_189 ;
wire \top/processor/sha_core/n3512_191 ;
wire \top/processor/sha_core/n3513_189 ;
wire \top/processor/sha_core/n3513_191 ;
wire \top/processor/sha_core/n3514_189 ;
wire \top/processor/sha_core/n3514_191 ;
wire \top/processor/sha_core/n3515_189 ;
wire \top/processor/sha_core/n3515_191 ;
wire \top/processor/sha_core/n3516_189 ;
wire \top/processor/sha_core/n3516_191 ;
wire \top/processor/sha_core/n3517_189 ;
wire \top/processor/sha_core/n3517_191 ;
wire \top/processor/sha_core/n3518_189 ;
wire \top/processor/sha_core/n3518_191 ;
wire \top/processor/sha_core/n3519_189 ;
wire \top/processor/sha_core/n3519_191 ;
wire \top/processor/sha_core/n3860_141 ;
wire \top/processor/sha_core/n3860_143 ;
wire \top/processor/sha_core/n3861_141 ;
wire \top/processor/sha_core/n3861_143 ;
wire \top/processor/sha_core/n3862_141 ;
wire \top/processor/sha_core/n3862_143 ;
wire \top/processor/sha_core/n3863_141 ;
wire \top/processor/sha_core/n3863_143 ;
wire \top/processor/sha_core/n3864_141 ;
wire \top/processor/sha_core/n3864_143 ;
wire \top/processor/sha_core/n3865_141 ;
wire \top/processor/sha_core/n3865_143 ;
wire \top/processor/sha_core/n3866_141 ;
wire \top/processor/sha_core/n3866_143 ;
wire \top/processor/sha_core/n3867_141 ;
wire \top/processor/sha_core/n3867_143 ;
wire \top/processor/sha_core/n3868_141 ;
wire \top/processor/sha_core/n3868_143 ;
wire \top/processor/sha_core/n3869_141 ;
wire \top/processor/sha_core/n3869_143 ;
wire \top/processor/sha_core/n3870_141 ;
wire \top/processor/sha_core/n3870_143 ;
wire \top/processor/sha_core/n3871_141 ;
wire \top/processor/sha_core/n3871_143 ;
wire \top/processor/sha_core/n3872_141 ;
wire \top/processor/sha_core/n3872_143 ;
wire \top/processor/sha_core/n3873_141 ;
wire \top/processor/sha_core/n3873_143 ;
wire \top/processor/sha_core/n3874_141 ;
wire \top/processor/sha_core/n3874_143 ;
wire \top/processor/sha_core/n3875_141 ;
wire \top/processor/sha_core/n3875_143 ;
wire \top/processor/sha_core/n3876_141 ;
wire \top/processor/sha_core/n3876_143 ;
wire \top/processor/sha_core/n3877_141 ;
wire \top/processor/sha_core/n3877_143 ;
wire \top/processor/sha_core/n3878_141 ;
wire \top/processor/sha_core/n3878_143 ;
wire \top/processor/sha_core/n3879_141 ;
wire \top/processor/sha_core/n3879_143 ;
wire \top/processor/sha_core/n3880_141 ;
wire \top/processor/sha_core/n3880_143 ;
wire \top/processor/sha_core/n3881_141 ;
wire \top/processor/sha_core/n3881_143 ;
wire \top/processor/sha_core/n3882_141 ;
wire \top/processor/sha_core/n3882_143 ;
wire \top/processor/sha_core/n3883_141 ;
wire \top/processor/sha_core/n3883_143 ;
wire \top/processor/sha_core/n3884_141 ;
wire \top/processor/sha_core/n3884_143 ;
wire \top/processor/sha_core/n3885_141 ;
wire \top/processor/sha_core/n3885_143 ;
wire \top/processor/sha_core/n3886_141 ;
wire \top/processor/sha_core/n3886_143 ;
wire \top/processor/sha_core/n3887_141 ;
wire \top/processor/sha_core/n3887_143 ;
wire \top/processor/sha_core/n3888_141 ;
wire \top/processor/sha_core/n3888_143 ;
wire \top/processor/sha_core/n3889_141 ;
wire \top/processor/sha_core/n3889_143 ;
wire \top/processor/sha_core/n3890_141 ;
wire \top/processor/sha_core/n3890_143 ;
wire \top/processor/sha_core/n3891_141 ;
wire \top/processor/sha_core/n3891_143 ;
wire \top/processor/sha_core/n327_213 ;
wire \top/processor/sha_core/n327_215 ;
wire \top/processor/sha_core/n327_217 ;
wire \top/processor/sha_core/n327_219 ;
wire \top/processor/sha_core/n328_213 ;
wire \top/processor/sha_core/n328_215 ;
wire \top/processor/sha_core/n328_217 ;
wire \top/processor/sha_core/n328_219 ;
wire \top/processor/sha_core/n329_213 ;
wire \top/processor/sha_core/n329_215 ;
wire \top/processor/sha_core/n329_217 ;
wire \top/processor/sha_core/n329_219 ;
wire \top/processor/sha_core/n330_213 ;
wire \top/processor/sha_core/n330_215 ;
wire \top/processor/sha_core/n330_217 ;
wire \top/processor/sha_core/n330_219 ;
wire \top/processor/sha_core/n331_213 ;
wire \top/processor/sha_core/n331_215 ;
wire \top/processor/sha_core/n331_217 ;
wire \top/processor/sha_core/n331_219 ;
wire \top/processor/sha_core/n332_213 ;
wire \top/processor/sha_core/n332_215 ;
wire \top/processor/sha_core/n332_217 ;
wire \top/processor/sha_core/n332_219 ;
wire \top/processor/sha_core/n333_213 ;
wire \top/processor/sha_core/n333_215 ;
wire \top/processor/sha_core/n333_217 ;
wire \top/processor/sha_core/n333_219 ;
wire \top/processor/sha_core/n334_213 ;
wire \top/processor/sha_core/n334_215 ;
wire \top/processor/sha_core/n334_217 ;
wire \top/processor/sha_core/n334_219 ;
wire \top/processor/sha_core/n335_213 ;
wire \top/processor/sha_core/n335_215 ;
wire \top/processor/sha_core/n335_217 ;
wire \top/processor/sha_core/n335_219 ;
wire \top/processor/sha_core/n336_213 ;
wire \top/processor/sha_core/n336_215 ;
wire \top/processor/sha_core/n336_217 ;
wire \top/processor/sha_core/n336_219 ;
wire \top/processor/sha_core/n337_213 ;
wire \top/processor/sha_core/n337_215 ;
wire \top/processor/sha_core/n337_217 ;
wire \top/processor/sha_core/n337_219 ;
wire \top/processor/sha_core/n338_213 ;
wire \top/processor/sha_core/n338_215 ;
wire \top/processor/sha_core/n338_217 ;
wire \top/processor/sha_core/n338_219 ;
wire \top/processor/sha_core/n339_213 ;
wire \top/processor/sha_core/n339_215 ;
wire \top/processor/sha_core/n339_217 ;
wire \top/processor/sha_core/n339_219 ;
wire \top/processor/sha_core/n340_213 ;
wire \top/processor/sha_core/n340_215 ;
wire \top/processor/sha_core/n340_217 ;
wire \top/processor/sha_core/n340_219 ;
wire \top/processor/sha_core/n341_213 ;
wire \top/processor/sha_core/n341_215 ;
wire \top/processor/sha_core/n341_217 ;
wire \top/processor/sha_core/n341_219 ;
wire \top/processor/sha_core/n342_213 ;
wire \top/processor/sha_core/n342_215 ;
wire \top/processor/sha_core/n342_217 ;
wire \top/processor/sha_core/n342_219 ;
wire \top/processor/sha_core/n343_213 ;
wire \top/processor/sha_core/n343_215 ;
wire \top/processor/sha_core/n343_217 ;
wire \top/processor/sha_core/n343_219 ;
wire \top/processor/sha_core/n344_213 ;
wire \top/processor/sha_core/n344_215 ;
wire \top/processor/sha_core/n344_217 ;
wire \top/processor/sha_core/n344_219 ;
wire \top/processor/sha_core/n345_213 ;
wire \top/processor/sha_core/n345_215 ;
wire \top/processor/sha_core/n345_217 ;
wire \top/processor/sha_core/n345_219 ;
wire \top/processor/sha_core/n346_213 ;
wire \top/processor/sha_core/n346_215 ;
wire \top/processor/sha_core/n346_217 ;
wire \top/processor/sha_core/n346_219 ;
wire \top/processor/sha_core/n347_213 ;
wire \top/processor/sha_core/n347_215 ;
wire \top/processor/sha_core/n347_217 ;
wire \top/processor/sha_core/n347_219 ;
wire \top/processor/sha_core/n348_213 ;
wire \top/processor/sha_core/n348_215 ;
wire \top/processor/sha_core/n348_217 ;
wire \top/processor/sha_core/n348_219 ;
wire \top/processor/sha_core/n349_213 ;
wire \top/processor/sha_core/n349_215 ;
wire \top/processor/sha_core/n349_217 ;
wire \top/processor/sha_core/n349_219 ;
wire \top/processor/sha_core/n350_213 ;
wire \top/processor/sha_core/n350_215 ;
wire \top/processor/sha_core/n350_217 ;
wire \top/processor/sha_core/n350_219 ;
wire \top/processor/sha_core/n351_213 ;
wire \top/processor/sha_core/n351_215 ;
wire \top/processor/sha_core/n351_217 ;
wire \top/processor/sha_core/n351_219 ;
wire \top/processor/sha_core/n352_213 ;
wire \top/processor/sha_core/n352_215 ;
wire \top/processor/sha_core/n352_217 ;
wire \top/processor/sha_core/n352_219 ;
wire \top/processor/sha_core/n353_213 ;
wire \top/processor/sha_core/n353_215 ;
wire \top/processor/sha_core/n353_217 ;
wire \top/processor/sha_core/n353_219 ;
wire \top/processor/sha_core/n354_213 ;
wire \top/processor/sha_core/n354_215 ;
wire \top/processor/sha_core/n354_217 ;
wire \top/processor/sha_core/n354_219 ;
wire \top/processor/sha_core/n355_213 ;
wire \top/processor/sha_core/n355_215 ;
wire \top/processor/sha_core/n355_217 ;
wire \top/processor/sha_core/n355_219 ;
wire \top/processor/sha_core/n356_213 ;
wire \top/processor/sha_core/n356_215 ;
wire \top/processor/sha_core/n356_217 ;
wire \top/processor/sha_core/n356_219 ;
wire \top/processor/sha_core/n357_213 ;
wire \top/processor/sha_core/n357_215 ;
wire \top/processor/sha_core/n357_217 ;
wire \top/processor/sha_core/n357_219 ;
wire \top/processor/sha_core/n358_213 ;
wire \top/processor/sha_core/n358_215 ;
wire \top/processor/sha_core/n358_217 ;
wire \top/processor/sha_core/n358_219 ;
wire \top/processor/sha_core/n3488_193 ;
wire \top/processor/sha_core/n3489_193 ;
wire \top/processor/sha_core/n3490_193 ;
wire \top/processor/sha_core/n3491_193 ;
wire \top/processor/sha_core/n3492_193 ;
wire \top/processor/sha_core/n3493_193 ;
wire \top/processor/sha_core/n3494_194 ;
wire \top/processor/sha_core/n3495_193 ;
wire \top/processor/sha_core/n3496_193 ;
wire \top/processor/sha_core/n3497_193 ;
wire \top/processor/sha_core/n3498_193 ;
wire \top/processor/sha_core/n3499_193 ;
wire \top/processor/sha_core/n3500_193 ;
wire \top/processor/sha_core/n3501_193 ;
wire \top/processor/sha_core/n3502_193 ;
wire \top/processor/sha_core/n3503_193 ;
wire \top/processor/sha_core/n3504_193 ;
wire \top/processor/sha_core/n3505_193 ;
wire \top/processor/sha_core/n3506_193 ;
wire \top/processor/sha_core/n3507_193 ;
wire \top/processor/sha_core/n3508_193 ;
wire \top/processor/sha_core/n3509_193 ;
wire \top/processor/sha_core/n3511_193 ;
wire \top/processor/sha_core/n3512_193 ;
wire \top/processor/sha_core/n3513_193 ;
wire \top/processor/sha_core/n3514_193 ;
wire \top/processor/sha_core/n3515_193 ;
wire \top/processor/sha_core/n3516_193 ;
wire \top/processor/sha_core/n3517_193 ;
wire \top/processor/sha_core/n3518_193 ;
wire \top/processor/sha_core/n3519_193 ;
wire \top/processor/sha_core/n3860_145 ;
wire \top/processor/sha_core/n3861_145 ;
wire \top/processor/sha_core/n3862_145 ;
wire \top/processor/sha_core/n3863_145 ;
wire \top/processor/sha_core/n3864_145 ;
wire \top/processor/sha_core/n3865_145 ;
wire \top/processor/sha_core/n3866_145 ;
wire \top/processor/sha_core/n3867_145 ;
wire \top/processor/sha_core/n3868_145 ;
wire \top/processor/sha_core/n3869_145 ;
wire \top/processor/sha_core/n3870_145 ;
wire \top/processor/sha_core/n3871_145 ;
wire \top/processor/sha_core/n3872_145 ;
wire \top/processor/sha_core/n3873_145 ;
wire \top/processor/sha_core/n3874_145 ;
wire \top/processor/sha_core/n3875_145 ;
wire \top/processor/sha_core/n3876_145 ;
wire \top/processor/sha_core/n3877_145 ;
wire \top/processor/sha_core/n3878_145 ;
wire \top/processor/sha_core/n3879_145 ;
wire \top/processor/sha_core/n3880_145 ;
wire \top/processor/sha_core/n3881_145 ;
wire \top/processor/sha_core/n3882_145 ;
wire \top/processor/sha_core/n3883_145 ;
wire \top/processor/sha_core/n3884_145 ;
wire \top/processor/sha_core/n3885_145 ;
wire \top/processor/sha_core/n3886_145 ;
wire \top/processor/sha_core/n3887_145 ;
wire \top/processor/sha_core/n3888_145 ;
wire \top/processor/sha_core/n3889_145 ;
wire \top/processor/sha_core/n3890_145 ;
wire \top/processor/sha_core/n3891_145 ;
wire \top/processor/sha_core/n327_221 ;
wire \top/processor/sha_core/n327_223 ;
wire \top/processor/sha_core/n328_221 ;
wire \top/processor/sha_core/n328_223 ;
wire \top/processor/sha_core/n329_221 ;
wire \top/processor/sha_core/n329_223 ;
wire \top/processor/sha_core/n330_221 ;
wire \top/processor/sha_core/n330_223 ;
wire \top/processor/sha_core/n331_221 ;
wire \top/processor/sha_core/n331_223 ;
wire \top/processor/sha_core/n332_221 ;
wire \top/processor/sha_core/n332_223 ;
wire \top/processor/sha_core/n333_221 ;
wire \top/processor/sha_core/n333_223 ;
wire \top/processor/sha_core/n334_221 ;
wire \top/processor/sha_core/n334_223 ;
wire \top/processor/sha_core/n335_221 ;
wire \top/processor/sha_core/n335_223 ;
wire \top/processor/sha_core/n336_221 ;
wire \top/processor/sha_core/n336_223 ;
wire \top/processor/sha_core/n337_221 ;
wire \top/processor/sha_core/n337_223 ;
wire \top/processor/sha_core/n338_221 ;
wire \top/processor/sha_core/n338_223 ;
wire \top/processor/sha_core/n339_221 ;
wire \top/processor/sha_core/n339_223 ;
wire \top/processor/sha_core/n340_221 ;
wire \top/processor/sha_core/n340_223 ;
wire \top/processor/sha_core/n341_221 ;
wire \top/processor/sha_core/n341_223 ;
wire \top/processor/sha_core/n342_221 ;
wire \top/processor/sha_core/n342_223 ;
wire \top/processor/sha_core/n343_221 ;
wire \top/processor/sha_core/n343_223 ;
wire \top/processor/sha_core/n344_221 ;
wire \top/processor/sha_core/n344_223 ;
wire \top/processor/sha_core/n345_221 ;
wire \top/processor/sha_core/n345_223 ;
wire \top/processor/sha_core/n346_221 ;
wire \top/processor/sha_core/n346_223 ;
wire \top/processor/sha_core/n347_221 ;
wire \top/processor/sha_core/n347_223 ;
wire \top/processor/sha_core/n348_221 ;
wire \top/processor/sha_core/n348_223 ;
wire \top/processor/sha_core/n349_221 ;
wire \top/processor/sha_core/n349_223 ;
wire \top/processor/sha_core/n350_221 ;
wire \top/processor/sha_core/n350_223 ;
wire \top/processor/sha_core/n351_221 ;
wire \top/processor/sha_core/n351_223 ;
wire \top/processor/sha_core/n352_221 ;
wire \top/processor/sha_core/n352_223 ;
wire \top/processor/sha_core/n353_221 ;
wire \top/processor/sha_core/n353_223 ;
wire \top/processor/sha_core/n354_221 ;
wire \top/processor/sha_core/n354_223 ;
wire \top/processor/sha_core/n355_221 ;
wire \top/processor/sha_core/n355_223 ;
wire \top/processor/sha_core/n356_221 ;
wire \top/processor/sha_core/n356_223 ;
wire \top/processor/sha_core/n357_221 ;
wire \top/processor/sha_core/n357_223 ;
wire \top/processor/sha_core/n358_221 ;
wire \top/processor/sha_core/n358_223 ;
wire \top/processor/sha_core/n3607_181 ;
wire \top/processor/sha_core/n3607_183 ;
wire \top/processor/sha_core/n3607_185 ;
wire \top/processor/sha_core/n3608_181 ;
wire \top/processor/sha_core/n3608_183 ;
wire \top/processor/sha_core/n3608_185 ;
wire \top/processor/sha_core/n3609_181 ;
wire \top/processor/sha_core/n3609_183 ;
wire \top/processor/sha_core/n3609_185 ;
wire \top/processor/sha_core/n3610_181 ;
wire \top/processor/sha_core/n3610_183 ;
wire \top/processor/sha_core/n3610_185 ;
wire \top/processor/sha_core/n3611_181 ;
wire \top/processor/sha_core/n3611_183 ;
wire \top/processor/sha_core/n3611_185 ;
wire \top/processor/sha_core/n3612_181 ;
wire \top/processor/sha_core/n3612_183 ;
wire \top/processor/sha_core/n3612_185 ;
wire \top/processor/sha_core/n3613_181 ;
wire \top/processor/sha_core/n3613_183 ;
wire \top/processor/sha_core/n3613_185 ;
wire \top/processor/sha_core/n3614_181 ;
wire \top/processor/sha_core/n3614_183 ;
wire \top/processor/sha_core/n3614_185 ;
wire \top/processor/sha_core/n3615_181 ;
wire \top/processor/sha_core/n3615_183 ;
wire \top/processor/sha_core/n3615_185 ;
wire \top/processor/sha_core/n3616_181 ;
wire \top/processor/sha_core/n3616_183 ;
wire \top/processor/sha_core/n3616_185 ;
wire \top/processor/sha_core/n3617_181 ;
wire \top/processor/sha_core/n3617_183 ;
wire \top/processor/sha_core/n3617_185 ;
wire \top/processor/sha_core/n3618_181 ;
wire \top/processor/sha_core/n3618_183 ;
wire \top/processor/sha_core/n3618_185 ;
wire \top/processor/sha_core/n3619_181 ;
wire \top/processor/sha_core/n3619_183 ;
wire \top/processor/sha_core/n3619_185 ;
wire \top/processor/sha_core/n3620_181 ;
wire \top/processor/sha_core/n3620_183 ;
wire \top/processor/sha_core/n3620_185 ;
wire \top/processor/sha_core/n3621_181 ;
wire \top/processor/sha_core/n3621_183 ;
wire \top/processor/sha_core/n3621_185 ;
wire \top/processor/sha_core/n3622_181 ;
wire \top/processor/sha_core/n3622_183 ;
wire \top/processor/sha_core/n3622_185 ;
wire \top/processor/sha_core/n3623_181 ;
wire \top/processor/sha_core/n3623_183 ;
wire \top/processor/sha_core/n3623_185 ;
wire \top/processor/sha_core/n3624_181 ;
wire \top/processor/sha_core/n3624_183 ;
wire \top/processor/sha_core/n3624_185 ;
wire \top/processor/sha_core/n3625_181 ;
wire \top/processor/sha_core/n3625_183 ;
wire \top/processor/sha_core/n3625_185 ;
wire \top/processor/sha_core/n3626_181 ;
wire \top/processor/sha_core/n3626_183 ;
wire \top/processor/sha_core/n3626_185 ;
wire \top/processor/sha_core/n3627_181 ;
wire \top/processor/sha_core/n3627_183 ;
wire \top/processor/sha_core/n3627_185 ;
wire \top/processor/sha_core/n3628_181 ;
wire \top/processor/sha_core/n3628_183 ;
wire \top/processor/sha_core/n3628_185 ;
wire \top/processor/sha_core/n3629_181 ;
wire \top/processor/sha_core/n3629_183 ;
wire \top/processor/sha_core/n3629_185 ;
wire \top/processor/sha_core/n3630_181 ;
wire \top/processor/sha_core/n3630_183 ;
wire \top/processor/sha_core/n3630_185 ;
wire \top/processor/sha_core/n3631_181 ;
wire \top/processor/sha_core/n3631_183 ;
wire \top/processor/sha_core/n3631_185 ;
wire \top/processor/sha_core/n3632_181 ;
wire \top/processor/sha_core/n3632_183 ;
wire \top/processor/sha_core/n3632_185 ;
wire \top/processor/sha_core/n3633_181 ;
wire \top/processor/sha_core/n3633_183 ;
wire \top/processor/sha_core/n3633_185 ;
wire \top/processor/sha_core/n3634_181 ;
wire \top/processor/sha_core/n3634_183 ;
wire \top/processor/sha_core/n3634_185 ;
wire \top/processor/sha_core/n3635_181 ;
wire \top/processor/sha_core/n3635_183 ;
wire \top/processor/sha_core/n3635_185 ;
wire \top/processor/sha_core/n3636_181 ;
wire \top/processor/sha_core/n3636_183 ;
wire \top/processor/sha_core/n3636_185 ;
wire \top/processor/sha_core/n3637_181 ;
wire \top/processor/sha_core/n3637_183 ;
wire \top/processor/sha_core/n3637_185 ;
wire \top/processor/sha_core/n3638_181 ;
wire \top/processor/sha_core/n3638_183 ;
wire \top/processor/sha_core/n3638_185 ;
wire [6:0] \top/processor/sha_core/msg_idx ;
wire [31:0] \top/processor/sha_core/w[0] ;
wire [31:0] \top/processor/sha_core/w[1] ;
wire [31:0] \top/processor/sha_core/w[2] ;
wire [31:0] \top/processor/sha_core/w[3] ;
wire [31:0] \top/processor/sha_core/w[4] ;
wire [31:0] \top/processor/sha_core/w[5] ;
wire [31:0] \top/processor/sha_core/w[6] ;
wire [31:0] \top/processor/sha_core/w[7] ;
wire [31:0] \top/processor/sha_core/w[8] ;
wire [31:0] \top/processor/sha_core/w[9] ;
wire [31:0] \top/processor/sha_core/w[10] ;
wire [31:0] \top/processor/sha_core/w[11] ;
wire [31:0] \top/processor/sha_core/w[12] ;
wire [31:0] \top/processor/sha_core/w[13] ;
wire [31:0] \top/processor/sha_core/w[14] ;
wire [31:0] \top/processor/sha_core/w[15] ;
wire [31:0] \top/processor/sha_core/w[16] ;
wire [31:0] \top/processor/sha_core/w[17] ;
wire [31:0] \top/processor/sha_core/w[18] ;
wire [31:0] \top/processor/sha_core/w[19] ;
wire [31:0] \top/processor/sha_core/w[20] ;
wire [31:0] \top/processor/sha_core/w[21] ;
wire [31:0] \top/processor/sha_core/w[22] ;
wire [31:0] \top/processor/sha_core/w[23] ;
wire [31:0] \top/processor/sha_core/w[24] ;
wire [31:0] \top/processor/sha_core/w[25] ;
wire [31:0] \top/processor/sha_core/w[26] ;
wire [31:0] \top/processor/sha_core/w[27] ;
wire [31:0] \top/processor/sha_core/w[28] ;
wire [31:0] \top/processor/sha_core/w[29] ;
wire [31:0] \top/processor/sha_core/w[30] ;
wire [31:0] \top/processor/sha_core/w[31] ;
wire [31:0] \top/processor/sha_core/w[32] ;
wire [31:0] \top/processor/sha_core/w[33] ;
wire [31:0] \top/processor/sha_core/w[34] ;
wire [31:0] \top/processor/sha_core/w[35] ;
wire [31:0] \top/processor/sha_core/w[36] ;
wire [31:0] \top/processor/sha_core/w[37] ;
wire [31:0] \top/processor/sha_core/w[38] ;
wire [31:0] \top/processor/sha_core/w[39] ;
wire [31:0] \top/processor/sha_core/w[40] ;
wire [31:0] \top/processor/sha_core/w[41] ;
wire [31:0] \top/processor/sha_core/w[42] ;
wire [31:0] \top/processor/sha_core/w[43] ;
wire [31:0] \top/processor/sha_core/w[44] ;
wire [31:0] \top/processor/sha_core/w[45] ;
wire [31:0] \top/processor/sha_core/w[46] ;
wire [31:0] \top/processor/sha_core/w[47] ;
wire [31:0] \top/processor/sha_core/w[48] ;
wire [31:0] \top/processor/sha_core/w[49] ;
wire [31:0] \top/processor/sha_core/w[50] ;
wire [31:0] \top/processor/sha_core/w[51] ;
wire [31:0] \top/processor/sha_core/w[52] ;
wire [31:0] \top/processor/sha_core/w[53] ;
wire [31:0] \top/processor/sha_core/w[54] ;
wire [31:0] \top/processor/sha_core/w[55] ;
wire [31:0] \top/processor/sha_core/w[56] ;
wire [31:0] \top/processor/sha_core/w[57] ;
wire [31:0] \top/processor/sha_core/w[58] ;
wire [31:0] \top/processor/sha_core/w[59] ;
wire [31:0] \top/processor/sha_core/w[60] ;
wire [31:0] \top/processor/sha_core/w[61] ;
wire [31:0] \top/processor/sha_core/w[62] ;
wire [31:0] \top/processor/sha_core/w[63] ;
wire [31:0] \top/processor/sha_core/h ;
wire [31:0] \top/processor/sha_core/g ;
wire [31:0] \top/processor/sha_core/f ;
wire [31:0] \top/processor/sha_core/e ;
wire [31:0] \top/processor/sha_core/d ;
wire [31:0] \top/processor/sha_core/c ;
wire [31:0] \top/processor/sha_core/b ;
wire [31:0] \top/processor/sha_core/a ;
wire [6:0] \top/processor/sha_core/t ;
wire [31:0] \top/processor/sha_core/h0 ;
wire [31:0] \top/processor/sha_core/h1 ;
wire [31:0] \top/processor/sha_core/h2 ;
wire [31:0] \top/processor/sha_core/h3 ;
wire [31:0] \top/processor/sha_core/h4 ;
wire [31:0] \top/processor/sha_core/h5 ;
wire [31:0] \top/processor/sha_core/h6 ;
wire [31:0] \top/processor/sha_core/h7 ;
wire [1:0] \top/processor/sha_core/state ;
VCC VCC_cZ (
  .V(VCC)
);
GND GND_cZ (
  .G(GND)
);
GSR GSR (
	.GSRI(VCC)
);
OBUF gowin_buf_0 (
	.I(uart_tx),
	.O(led0)
);
LUT3 \top/n568_s15  (
	.I0(\top/state [2]),
	.I1(\top/state [0]),
	.I2(\top/state [1]),
	.F(\top/n568_23 )
);
defparam \top/n568_s15 .INIT=8'hB4;
LUT2 \top/n635_s2  (
	.I0(rst),
	.I1(\top/n570_11 ),
	.F(\top/tx_data_4_15 )
);
defparam \top/n635_s2 .INIT=4'h4;
LUT3 \top/n636_s2  (
	.I0(\top/n523_6 ),
	.I1(\top/n523_5 ),
	.I2(\top/n522_5 ),
	.F(\top/n636_5 )
);
defparam \top/n636_s2 .INIT=8'h07;
LUT2 \top/data_in_7_s2  (
	.I0(rst),
	.I1(\top/n586_12 ),
	.F(\top/data_in_7_6 )
);
defparam \top/data_in_7_s2 .INIT=4'h4;
LUT4 \top/send_index_6_s3  (
	.I0(\top/state [2]),
	.I1(\top/state [1]),
	.I2(\top/send_index_6_8 ),
	.I3(\top/n570_11 ),
	.F(\top/send_index_6_7 )
);
defparam \top/send_index_6_s3 .INIT=16'hFF40;
LUT4 \top/n568_s16  (
	.I0(\top/n568_26 ),
	.I1(\top/n568_27 ),
	.I2(\top/n586_10 ),
	.I3(\top/n568_28 ),
	.F(\top/n568_25 )
);
defparam \top/n568_s16 .INIT=16'h00EF;
LUT2 \top/n585_s10  (
	.I0(\top/send_index [0]),
	.I1(\top/state [0]),
	.F(\top/n585_15 )
);
defparam \top/n585_s10 .INIT=4'h4;
LUT3 \top/n584_s9  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/state [0]),
	.F(\top/n584_14 )
);
defparam \top/n584_s9 .INIT=8'h60;
LUT3 \top/n582_s9  (
	.I0(\top/send_index [3]),
	.I1(\top/n582_17 ),
	.I2(\top/state [0]),
	.F(\top/n582_14 )
);
defparam \top/n582_s9 .INIT=8'h60;
LUT4 \top/n581_s9  (
	.I0(\top/send_index [3]),
	.I1(\top/n582_17 ),
	.I2(\top/send_index [4]),
	.I3(\top/state [0]),
	.F(\top/n581_14 )
);
defparam \top/n581_s9 .INIT=16'h7800;
LUT3 \top/n580_s9  (
	.I0(\top/send_index [5]),
	.I1(\top/n580_15 ),
	.I2(\top/state [0]),
	.F(\top/n580_14 )
);
defparam \top/n580_s9 .INIT=8'h60;
LUT4 \top/n579_s10  (
	.I0(\top/send_index [5]),
	.I1(\top/n580_15 ),
	.I2(\top/send_index [6]),
	.I3(\top/state [0]),
	.F(\top/n579_15 )
);
defparam \top/n579_s10 .INIT=16'h7800;
LUT3 \top/n567_s13  (
	.I0(\top/state [2]),
	.I1(\top/state [1]),
	.I2(\top/state [0]),
	.F(\top/n567_20 )
);
defparam \top/n567_s13 .INIT=8'h40;
LUT4 \top/n522_s1  (
	.I0(\top/n522_6 ),
	.I1(\top/n522_7 ),
	.I2(\top/n522_8 ),
	.I3(\top/n522_9 ),
	.F(\top/n522_5 )
);
defparam \top/n522_s1 .INIT=16'h8000;
LUT4 \top/n523_s2  (
	.I0(\top/n523_7 ),
	.I1(\top/n523_8 ),
	.I2(\top/n523_9 ),
	.I3(\top/n523_10 ),
	.F(\top/n523_5 )
);
defparam \top/n523_s2 .INIT=16'h8000;
LUT4 \top/n523_s3  (
	.I0(\top/n523_11 ),
	.I1(\top/n523_12 ),
	.I2(\top/n523_13 ),
	.I3(\top/n523_14 ),
	.F(\top/n523_6 )
);
defparam \top/n523_s3 .INIT=16'h8000;
LUT4 \top/n525_s1  (
	.I0(\top/n525_5 ),
	.I1(\top/n525_6 ),
	.I2(\top/n525_7 ),
	.I3(\top/n525_8 ),
	.F(\top/n525_4 )
);
defparam \top/n525_s1 .INIT=16'h8000;
LUT2 \top/n586_s6  (
	.I0(\top/state [1]),
	.I1(\top/state [2]),
	.F(\top/n586_10 )
);
defparam \top/n586_s6 .INIT=4'h1;
LUT3 \top/state_0_s4  (
	.I0(\top/state [0]),
	.I1(\top/state [1]),
	.I2(\top/tx_busy_Z ),
	.F(\top/state_0_9 )
);
defparam \top/state_0_s4 .INIT=8'h01;
LUT4 \top/send_index_6_s4  (
	.I0(\top/state [0]),
	.I1(\top/state_0 [0]),
	.I2(\top/state_0 [1]),
	.I3(\top/state_0 [2]),
	.F(\top/send_index_6_8 )
);
defparam \top/send_index_6_s4 .INIT=16'h0100;
LUT4 \top/n568_s17  (
	.I0(\top/n568_29 ),
	.I1(\top/rx_data_Z [0]),
	.I2(\top/rx_data_Z [1]),
	.I3(\top/n568_30 ),
	.F(\top/n568_26 )
);
defparam \top/n568_s17 .INIT=16'h8000;
LUT4 \top/n568_s18  (
	.I0(\top/rx_data_Z [1]),
	.I1(\top/rx_data_Z [0]),
	.I2(\top/n568_31 ),
	.I3(\top/n568_32 ),
	.F(\top/n568_27 )
);
defparam \top/n568_s18 .INIT=16'h4000;
LUT4 \top/n568_s19  (
	.I0(\top/n568_33 ),
	.I1(\top/state [2]),
	.I2(\top/send_index_6_8 ),
	.I3(\top/state [1]),
	.F(\top/n568_28 )
);
defparam \top/n568_s19 .INIT=16'h0100;
LUT2 \top/n583_s10  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.F(\top/n583_15 )
);
defparam \top/n583_s10 .INIT=4'h8;
LUT3 \top/n580_s10  (
	.I0(\top/send_index [3]),
	.I1(\top/send_index [4]),
	.I2(\top/n582_17 ),
	.F(\top/n580_15 )
);
defparam \top/n580_s10 .INIT=8'h80;
LUT4 \top/n522_s2  (
	.I0(\top/n522_10 ),
	.I1(\top/n522_11 ),
	.I2(\top/n522_12 ),
	.I3(\top/n522_13 ),
	.F(\top/n522_6 )
);
defparam \top/n522_s2 .INIT=16'h4000;
LUT4 \top/n522_s3  (
	.I0(\top/n522_14 ),
	.I1(\top/n522_94 ),
	.I2(\top/n522_16 ),
	.I3(\top/n522_17 ),
	.F(\top/n522_7 )
);
defparam \top/n522_s3 .INIT=16'h1000;
LUT4 \top/n522_s4  (
	.I0(\top/n522_18 ),
	.I1(\top/n522_19 ),
	.I2(\top/n522_20 ),
	.I3(\top/n522_21 ),
	.F(\top/n522_8 )
);
defparam \top/n522_s4 .INIT=16'h8000;
LUT4 \top/n522_s5  (
	.I0(\top/n522_22 ),
	.I1(\top/n522_23 ),
	.I2(\top/n522_24 ),
	.I3(\top/n522_25 ),
	.F(\top/n522_9 )
);
defparam \top/n522_s5 .INIT=16'h4000;
LUT4 \top/n523_s4  (
	.I0(\top/n523_15 ),
	.I1(\top/n523_16 ),
	.I2(\top/n523_17 ),
	.I3(\top/n523_18 ),
	.F(\top/n523_7 )
);
defparam \top/n523_s4 .INIT=16'h4000;
LUT4 \top/n523_s5  (
	.I0(\top/n523_19 ),
	.I1(\top/n523_20 ),
	.I2(\top/n523_21 ),
	.I3(\top/n523_22 ),
	.F(\top/n523_8 )
);
defparam \top/n523_s5 .INIT=16'h8000;
LUT4 \top/n523_s6  (
	.I0(\top/n523_23 ),
	.I1(\top/n523_24 ),
	.I2(\top/n523_25 ),
	.I3(\top/n523_26 ),
	.F(\top/n523_9 )
);
defparam \top/n523_s6 .INIT=16'h1000;
LUT4 \top/n523_s7  (
	.I0(\top/n523_27 ),
	.I1(\top/n523_28 ),
	.I2(\top/n523_29 ),
	.I3(\top/n523_30 ),
	.F(\top/n523_10 )
);
defparam \top/n523_s7 .INIT=16'h4000;
LUT4 \top/n523_s8  (
	.I0(\top/n523_31 ),
	.I1(\top/n523_32 ),
	.I2(\top/n523_33 ),
	.I3(\top/n523_34 ),
	.F(\top/n523_11 )
);
defparam \top/n523_s8 .INIT=16'h8000;
LUT4 \top/n523_s9  (
	.I0(\top/n523_35 ),
	.I1(\top/n523_36 ),
	.I2(\top/n523_37 ),
	.I3(\top/n523_38 ),
	.F(\top/n523_12 )
);
defparam \top/n523_s9 .INIT=16'h4000;
LUT4 \top/n523_s10  (
	.I0(\top/n523_39 ),
	.I1(\top/n523_40 ),
	.I2(\top/n523_41 ),
	.I3(\top/n523_42 ),
	.F(\top/n523_13 )
);
defparam \top/n523_s10 .INIT=16'h4000;
LUT4 \top/n523_s11  (
	.I0(\top/n523_43 ),
	.I1(\top/n523_44 ),
	.I2(\top/n523_45 ),
	.I3(\top/n523_46 ),
	.F(\top/n523_14 )
);
defparam \top/n523_s11 .INIT=16'h1000;
LUT4 \top/n525_s2  (
	.I0(\top/n525_9 ),
	.I1(\top/n525_10 ),
	.I2(\top/n525_11 ),
	.I3(\top/n525_12 ),
	.F(\top/n525_5 )
);
defparam \top/n525_s2 .INIT=16'h1000;
LUT4 \top/n525_s3  (
	.I0(\top/n525_13 ),
	.I1(\top/n525_14 ),
	.I2(\top/n525_15 ),
	.I3(\top/n525_16 ),
	.F(\top/n525_6 )
);
defparam \top/n525_s3 .INIT=16'h8000;
LUT4 \top/n525_s4  (
	.I0(\top/n525_17 ),
	.I1(\top/n525_18 ),
	.I2(\top/n525_19 ),
	.I3(\top/n525_20 ),
	.F(\top/n525_7 )
);
defparam \top/n525_s4 .INIT=16'h4000;
LUT4 \top/n525_s5  (
	.I0(\top/n525_21 ),
	.I1(\top/n525_22 ),
	.I2(\top/n525_23 ),
	.I3(\top/n525_24 ),
	.F(\top/n525_8 )
);
defparam \top/n525_s5 .INIT=16'h4000;
LUT4 \top/n568_s20  (
	.I0(\top/rx_data_Z [2]),
	.I1(\top/rx_data_Z [3]),
	.I2(\top/rx_data_Z [4]),
	.I3(\top/rx_data_Z [5]),
	.F(\top/n568_29 )
);
defparam \top/n568_s20 .INIT=16'h8000;
LUT4 \top/n568_s21  (
	.I0(\top/rx_data_Z [6]),
	.I1(\top/rx_data_Z [7]),
	.I2(\top/rx_valid_Z ),
	.I3(\top/state [0]),
	.F(\top/n568_30 )
);
defparam \top/n568_s21 .INIT=16'h8000;
LUT4 \top/n568_s22  (
	.I0(\top/rx_data_Z [2]),
	.I1(\top/rx_data_Z [3]),
	.I2(\top/rx_data_Z [4]),
	.I3(\top/rx_data_Z [5]),
	.F(\top/n568_31 )
);
defparam \top/n568_s22 .INIT=16'h0001;
LUT4 \top/n568_s23  (
	.I0(\top/rx_data_Z [6]),
	.I1(\top/rx_data_Z [7]),
	.I2(\top/state [0]),
	.I3(\top/rx_valid_Z ),
	.F(\top/n568_32 )
);
defparam \top/n568_s23 .INIT=16'h0100;
LUT4 \top/n568_s24  (
	.I0(\top/tx_busy_Z ),
	.I1(\top/state [0]),
	.I2(\top/n568_34 ),
	.I3(\top/n582_17 ),
	.F(\top/n568_33 )
);
defparam \top/n568_s24 .INIT=16'h4000;
LUT4 \top/n522_s6  (
	.I0(\top/n522_26 ),
	.I1(\top/n522_27 ),
	.I2(\top/n522_28 ),
	.I3(\top/n568_34 ),
	.F(\top/n522_10 )
);
defparam \top/n522_s6 .INIT=16'hF800;
LUT4 \top/n522_s7  (
	.I0(\top/n522_29 ),
	.I1(\top/n522_30 ),
	.I2(\top/n522_31 ),
	.I3(\top/n522_32 ),
	.F(\top/n522_11 )
);
defparam \top/n522_s7 .INIT=16'h008F;
LUT4 \top/n522_s8  (
	.I0(\top/n522_33 ),
	.I1(\top/n522_34 ),
	.I2(\top/n522_35 ),
	.I3(\top/n522_36 ),
	.F(\top/n522_12 )
);
defparam \top/n522_s8 .INIT=16'h0001;
LUT4 \top/n522_s9  (
	.I0(\top/n522_37 ),
	.I1(\top/n522_38 ),
	.I2(\top/n522_39 ),
	.I3(\top/n522_40 ),
	.F(\top/n522_13 )
);
defparam \top/n522_s9 .INIT=16'h000B;
LUT4 \top/n522_s10  (
	.I0(\top/n522_41 ),
	.I1(\top/n522_42 ),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n522_14 )
);
defparam \top/n522_s10 .INIT=16'h0C0A;
LUT4 \top/n522_s12  (
	.I0(\top/hash_out [39]),
	.I1(\top/n522_38 ),
	.I2(\top/n522_45 ),
	.I3(\top/n522_46 ),
	.F(\top/n522_16 )
);
defparam \top/n522_s12 .INIT=16'h007F;
LUT4 \top/n522_s13  (
	.I0(\top/send_index [2]),
	.I1(\top/n522_47 ),
	.I2(\top/n522_48 ),
	.I3(\top/n522_49 ),
	.F(\top/n522_17 )
);
defparam \top/n522_s13 .INIT=16'h00EF;
LUT4 \top/n522_s14  (
	.I0(\top/n522_50 ),
	.I1(\top/n522_51 ),
	.I2(\top/n522_52 ),
	.I3(\top/n522_53 ),
	.F(\top/n522_18 )
);
defparam \top/n522_s14 .INIT=16'h0BBB;
LUT4 \top/n522_s15  (
	.I0(\top/n522_45 ),
	.I1(\top/n522_54 ),
	.I2(\top/n522_92 ),
	.I3(\top/send_index [2]),
	.F(\top/n522_19 )
);
defparam \top/n522_s15 .INIT=16'h0F77;
LUT4 \top/n522_s16  (
	.I0(\top/hash_out [243]),
	.I1(\top/n522_56 ),
	.I2(\top/n522_31 ),
	.I3(\top/n522_57 ),
	.F(\top/n522_20 )
);
defparam \top/n522_s16 .INIT=16'h007F;
LUT4 \top/n522_s17  (
	.I0(\top/n522_90 ),
	.I1(\top/hash_out [155]),
	.I2(\top/n522_59 ),
	.I3(\top/n522_60 ),
	.F(\top/n522_21 )
);
defparam \top/n522_s17 .INIT=16'h0007;
LUT4 \top/n522_s18  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [159]),
	.I2(\top/n522_61 ),
	.I3(\top/n522_62 ),
	.F(\top/n522_22 )
);
defparam \top/n522_s18 .INIT=16'h4000;
LUT4 \top/n522_s19  (
	.I0(\top/n522_63 ),
	.I1(\top/n522_64 ),
	.I2(\top/n522_65 ),
	.I3(\top/n522_66 ),
	.F(\top/n522_23 )
);
defparam \top/n522_s19 .INIT=16'h001F;
LUT4 \top/n522_s20  (
	.I0(\top/n522_67 ),
	.I1(\top/n522_52 ),
	.I2(\top/n522_68 ),
	.I3(\top/n522_69 ),
	.F(\top/n522_24 )
);
defparam \top/n522_s20 .INIT=16'h000B;
LUT4 \top/n522_s21  (
	.I0(\top/n522_70 ),
	.I1(\top/n522_71 ),
	.I2(\top/n522_72 ),
	.I3(\top/n522_73 ),
	.F(\top/n522_25 )
);
defparam \top/n522_s21 .INIT=16'h0001;
LUT4 \top/n523_s12  (
	.I0(\top/n523_47 ),
	.I1(\top/n523_48 ),
	.I2(\top/send_index [2]),
	.I3(\top/n568_34 ),
	.F(\top/n523_15 )
);
defparam \top/n523_s12 .INIT=16'hC500;
LUT4 \top/n523_s13  (
	.I0(\top/n523_49 ),
	.I1(\top/n522_45 ),
	.I2(\top/n523_50 ),
	.I3(\top/n523_153 ),
	.F(\top/n523_16 )
);
defparam \top/n523_s13 .INIT=16'h000B;
LUT4 \top/n523_s14  (
	.I0(\top/n523_52 ),
	.I1(\top/n522_38 ),
	.I2(\top/n523_53 ),
	.I3(\top/n523_54 ),
	.F(\top/n523_17 )
);
defparam \top/n523_s14 .INIT=16'h000B;
LUT3 \top/n523_s15  (
	.I0(\top/n523_55 ),
	.I1(\top/n522_48 ),
	.I2(\top/n523_56 ),
	.F(\top/n523_18 )
);
defparam \top/n523_s15 .INIT=8'h0B;
LUT4 \top/n523_s16  (
	.I0(\top/n522_52 ),
	.I1(\top/n523_57 ),
	.I2(\top/n523_151 ),
	.I3(\top/send_index [2]),
	.F(\top/n523_19 )
);
defparam \top/n523_s16 .INIT=16'h770F;
LUT3 \top/n523_s17  (
	.I0(\top/n522_90 ),
	.I1(\top/hash_out [153]),
	.I2(\top/n523_59 ),
	.F(\top/n523_20 )
);
defparam \top/n523_s17 .INIT=8'h07;
LUT4 \top/n523_s18  (
	.I0(\top/n522_56 ),
	.I1(\top/n523_60 ),
	.I2(\top/n523_61 ),
	.I3(\top/n523_62 ),
	.F(\top/n523_21 )
);
defparam \top/n523_s18 .INIT=16'h000D;
LUT4 \top/n523_s19  (
	.I0(\top/hash_out [113]),
	.I1(\top/n522_65 ),
	.I2(\top/n522_31 ),
	.I3(\top/n523_63 ),
	.F(\top/n523_22 )
);
defparam \top/n523_s19 .INIT=16'h007F;
LUT4 \top/n523_s20  (
	.I0(\top/n523_64 ),
	.I1(\top/n523_65 ),
	.I2(\top/send_index [0]),
	.I3(\top/n522_56 ),
	.F(\top/n523_23 )
);
defparam \top/n523_s20 .INIT=16'h3500;
LUT4 \top/n523_s21  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [85]),
	.I2(\top/n523_66 ),
	.I3(\top/n522_52 ),
	.F(\top/n523_24 )
);
defparam \top/n523_s21 .INIT=16'h4000;
LUT2 \top/n523_s22  (
	.I0(\top/n523_67 ),
	.I1(\top/n523_68 ),
	.F(\top/n523_25 )
);
defparam \top/n523_s22 .INIT=4'h1;
LUT4 \top/n523_s23  (
	.I0(\top/n523_69 ),
	.I1(\top/n523_70 ),
	.I2(\top/n523_71 ),
	.I3(\top/n523_72 ),
	.F(\top/n523_26 )
);
defparam \top/n523_s23 .INIT=16'h0007;
LUT4 \top/n523_s24  (
	.I0(\top/n523_73 ),
	.I1(\top/send_index [0]),
	.I2(\top/n523_74 ),
	.I3(\top/send_index [2]),
	.F(\top/n523_27 )
);
defparam \top/n523_s24 .INIT=16'h0130;
LUT4 \top/n523_s25  (
	.I0(\top/n523_69 ),
	.I1(\top/n523_75 ),
	.I2(\top/n523_76 ),
	.I3(\top/n522_51 ),
	.F(\top/n523_28 )
);
defparam \top/n523_s25 .INIT=16'h0777;
LUT4 \top/n523_s26  (
	.I0(\top/n523_77 ),
	.I1(\top/n523_78 ),
	.I2(\top/n523_79 ),
	.I3(\top/n523_80 ),
	.F(\top/n523_29 )
);
defparam \top/n523_s26 .INIT=16'h000D;
LUT4 \top/n523_s27  (
	.I0(\top/n523_81 ),
	.I1(\top/n522_65 ),
	.I2(\top/send_index [2]),
	.I3(\top/n523_82 ),
	.F(\top/n523_30 )
);
defparam \top/n523_s27 .INIT=16'h00BF;
LUT4 \top/n523_s28  (
	.I0(\top/n523_83 ),
	.I1(\top/n523_84 ),
	.I2(\top/n523_85 ),
	.I3(\top/n523_86 ),
	.F(\top/n523_31 )
);
defparam \top/n523_s28 .INIT=16'h0100;
LUT4 \top/n523_s29  (
	.I0(\top/n523_87 ),
	.I1(\top/n523_88 ),
	.I2(\top/n523_89 ),
	.I3(\top/n523_90 ),
	.F(\top/n523_32 )
);
defparam \top/n523_s29 .INIT=16'h0007;
LUT4 \top/n523_s30  (
	.I0(\top/n523_91 ),
	.I1(\top/n522_51 ),
	.I2(\top/n523_92 ),
	.I3(\top/n523_93 ),
	.F(\top/n523_33 )
);
defparam \top/n523_s30 .INIT=16'h000B;
LUT4 \top/n523_s31  (
	.I0(\top/hash_out [118]),
	.I1(\top/n522_65 ),
	.I2(\top/n523_77 ),
	.I3(\top/n523_94 ),
	.F(\top/n523_34 )
);
defparam \top/n523_s31 .INIT=16'h007F;
LUT3 \top/n523_s32  (
	.I0(\top/n523_95 ),
	.I1(\top/n523_96 ),
	.I2(\top/n522_52 ),
	.F(\top/n523_35 )
);
defparam \top/n523_s32 .INIT=8'h70;
LUT4 \top/n523_s33  (
	.I0(\top/n523_97 ),
	.I1(\top/n523_88 ),
	.I2(\top/send_index [0]),
	.I3(\top/n523_98 ),
	.F(\top/n523_36 )
);
defparam \top/n523_s33 .INIT=16'h00BF;
LUT4 \top/n523_s34  (
	.I0(\top/n523_99 ),
	.I1(\top/n523_100 ),
	.I2(\top/n523_149 ),
	.I3(\top/n523_102 ),
	.F(\top/n523_37 )
);
defparam \top/n523_s34 .INIT=16'h0100;
LUT4 \top/n523_s35  (
	.I0(\top/n568_34 ),
	.I1(\top/n523_103 ),
	.I2(\top/send_index [2]),
	.I3(\top/n523_104 ),
	.F(\top/n523_38 )
);
defparam \top/n523_s35 .INIT=16'h00DF;
LUT4 \top/n523_s36  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [34]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_45 ),
	.F(\top/n523_39 )
);
defparam \top/n523_s36 .INIT=16'h8000;
LUT4 \top/n523_s37  (
	.I0(\top/n523_105 ),
	.I1(\top/n523_77 ),
	.I2(\top/n523_106 ),
	.I3(\top/n523_107 ),
	.F(\top/n523_40 )
);
defparam \top/n523_s37 .INIT=16'h000B;
LUT4 \top/n523_s38  (
	.I0(\top/hash_out [70]),
	.I1(\top/n522_38 ),
	.I2(\top/n522_52 ),
	.I3(\top/n523_108 ),
	.F(\top/n523_41 )
);
defparam \top/n523_s38 .INIT=16'h007F;
LUT4 \top/n523_s39  (
	.I0(\top/n523_109 ),
	.I1(\top/n523_110 ),
	.I2(\top/n523_111 ),
	.I3(\top/n523_112 ),
	.F(\top/n523_42 )
);
defparam \top/n523_s39 .INIT=16'h0001;
LUT4 \top/n523_s40  (
	.I0(\top/n523_113 ),
	.I1(\top/send_index [2]),
	.I2(\top/n523_114 ),
	.I3(\top/n522_45 ),
	.F(\top/n523_43 )
);
defparam \top/n523_s40 .INIT=16'h4F00;
LUT4 \top/n523_s41  (
	.I0(\top/n523_115 ),
	.I1(\top/n523_116 ),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n523_44 )
);
defparam \top/n523_s41 .INIT=16'h0A0C;
LUT4 \top/n523_s42  (
	.I0(\top/hash_out [142]),
	.I1(\top/n522_61 ),
	.I2(\top/n523_117 ),
	.I3(\top/n523_118 ),
	.F(\top/n523_45 )
);
defparam \top/n523_s42 .INIT=16'h007F;
LUT4 \top/n523_s43  (
	.I0(\top/n522_56 ),
	.I1(\top/n522_31 ),
	.I2(\top/hash_out [242]),
	.I3(\top/n523_119 ),
	.F(\top/n523_46 )
);
defparam \top/n523_s43 .INIT=16'h007F;
LUT4 \top/n525_s6  (
	.I0(\top/send_index [0]),
	.I1(\top/n525_25 ),
	.I2(\top/n525_26 ),
	.I3(\top/n522_51 ),
	.F(\top/n525_9 )
);
defparam \top/n525_s6 .INIT=16'hF800;
LUT4 \top/n525_s7  (
	.I0(\top/n525_27 ),
	.I1(\top/n525_28 ),
	.I2(\top/send_index [2]),
	.I3(\top/n568_34 ),
	.F(\top/n525_10 )
);
defparam \top/n525_s7 .INIT=16'h5C00;
LUT4 \top/n525_s8  (
	.I0(\top/n525_29 ),
	.I1(\top/n525_30 ),
	.I2(\top/n525_31 ),
	.I3(\top/n525_32 ),
	.F(\top/n525_11 )
);
defparam \top/n525_s8 .INIT=16'h0100;
LUT3 \top/n525_s9  (
	.I0(\top/n525_33 ),
	.I1(\top/n522_61 ),
	.I2(\top/n525_34 ),
	.F(\top/n525_12 )
);
defparam \top/n525_s9 .INIT=8'h07;
LUT3 \top/n525_s10  (
	.I0(\top/n525_35 ),
	.I1(\top/n522_56 ),
	.I2(\top/n525_36 ),
	.F(\top/n525_13 )
);
defparam \top/n525_s10 .INIT=8'h0B;
LUT4 \top/n525_s11  (
	.I0(\top/send_index [1]),
	.I1(\top/n525_37 ),
	.I2(\top/n522_61 ),
	.I3(\top/n525_38 ),
	.F(\top/n525_14 )
);
defparam \top/n525_s11 .INIT=16'hEF00;
LUT4 \top/n525_s12  (
	.I0(\top/n525_39 ),
	.I1(\top/n522_65 ),
	.I2(\top/send_index [0]),
	.I3(\top/n525_40 ),
	.F(\top/n525_15 )
);
defparam \top/n525_s12 .INIT=16'h00BF;
LUT4 \top/n525_s13  (
	.I0(\top/n525_41 ),
	.I1(\top/n522_44 ),
	.I2(\top/n525_42 ),
	.I3(\top/n525_43 ),
	.F(\top/n525_16 )
);
defparam \top/n525_s13 .INIT=16'h0007;
LUT4 \top/n525_s14  (
	.I0(\top/send_index [3]),
	.I1(\top/send_index [4]),
	.I2(\top/n525_44 ),
	.I3(\top/n522_31 ),
	.F(\top/n525_17 )
);
defparam \top/n525_s14 .INIT=16'h1000;
LUT4 \top/n525_s15  (
	.I0(\top/n525_45 ),
	.I1(\top/n522_51 ),
	.I2(\top/n525_46 ),
	.I3(\top/n525_47 ),
	.F(\top/n525_18 )
);
defparam \top/n525_s15 .INIT=16'h0007;
LUT2 \top/n525_s16  (
	.I0(\top/n525_48 ),
	.I1(\top/n525_49 ),
	.F(\top/n525_19 )
);
defparam \top/n525_s16 .INIT=4'h1;
LUT4 \top/n525_s17  (
	.I0(\top/n525_50 ),
	.I1(\top/n525_51 ),
	.I2(\top/n525_52 ),
	.I3(\top/n525_53 ),
	.F(\top/n525_20 )
);
defparam \top/n525_s17 .INIT=16'h000B;
LUT3 \top/n525_s18  (
	.I0(\top/n525_54 ),
	.I1(\top/n525_55 ),
	.I2(\top/n522_52 ),
	.F(\top/n525_21 )
);
defparam \top/n525_s18 .INIT=8'hB0;
LUT4 \top/n525_s19  (
	.I0(\top/n522_65 ),
	.I1(\top/n523_77 ),
	.I2(\top/hash_out [116]),
	.I3(\top/n525_56 ),
	.F(\top/n525_22 )
);
defparam \top/n525_s19 .INIT=16'h007F;
LUT3 \top/n525_s20  (
	.I0(\top/n525_57 ),
	.I1(\top/n522_31 ),
	.I2(\top/n525_58 ),
	.F(\top/n525_23 )
);
defparam \top/n525_s20 .INIT=8'h0B;
LUT4 \top/n525_s21  (
	.I0(\top/n525_59 ),
	.I1(\top/n523_77 ),
	.I2(\top/n525_60 ),
	.I3(\top/n525_61 ),
	.F(\top/n525_24 )
);
defparam \top/n525_s21 .INIT=16'h000B;
LUT4 \top/n568_s25  (
	.I0(\top/send_index [6]),
	.I1(\top/send_index [4]),
	.I2(\top/send_index [5]),
	.I3(\top/send_index [3]),
	.F(\top/n568_34 )
);
defparam \top/n568_s25 .INIT=16'h4000;
LUT4 \top/n522_s22  (
	.I0(\top/send_index [0]),
	.I1(\top/hash_out [31]),
	.I2(\top/n522_74 ),
	.I3(\top/send_index [1]),
	.F(\top/n522_26 )
);
defparam \top/n522_s22 .INIT=16'hF0EE;
LUT4 \top/n522_s23  (
	.I0(\top/send_index [1]),
	.I1(\top/hash_out [27]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [2]),
	.F(\top/n522_27 )
);
defparam \top/n522_s23 .INIT=16'h00EF;
LUT4 \top/n522_s24  (
	.I0(\top/send_index [0]),
	.I1(\top/hash_out [11]),
	.I2(\top/n522_75 ),
	.I3(\top/n522_76 ),
	.F(\top/n522_28 )
);
defparam \top/n522_s24 .INIT=16'hF800;
LUT4 \top/n522_s25  (
	.I0(\top/n522_48 ),
	.I1(\top/hash_out [211]),
	.I2(\top/hash_out [179]),
	.I3(\top/n522_51 ),
	.F(\top/n522_29 )
);
defparam \top/n522_s25 .INIT=16'h0777;
LUT4 \top/n522_s26  (
	.I0(\top/n522_61 ),
	.I1(\top/hash_out [147]),
	.I2(\top/n522_77 ),
	.I3(\top/n522_78 ),
	.F(\top/n522_30 )
);
defparam \top/n522_s26 .INIT=16'h0777;
LUT3 \top/n522_s27  (
	.I0(\top/send_index [2]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [0]),
	.F(\top/n522_31 )
);
defparam \top/n522_s27 .INIT=8'h40;
LUT4 \top/n522_s28  (
	.I0(\top/n522_79 ),
	.I1(\top/send_index [2]),
	.I2(\top/n522_80 ),
	.I3(\top/n583_15 ),
	.F(\top/n522_32 )
);
defparam \top/n522_s28 .INIT=16'h4000;
LUT3 \top/n522_s29  (
	.I0(\top/hash_out [71]),
	.I1(\top/n522_38 ),
	.I2(\top/n522_52 ),
	.F(\top/n522_33 )
);
defparam \top/n522_s29 .INIT=8'h80;
LUT4 \top/n522_s30  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [235]),
	.I2(\top/n522_56 ),
	.I3(\top/n522_44 ),
	.F(\top/n522_34 )
);
defparam \top/n522_s30 .INIT=16'h8000;
LUT4 \top/n522_s31  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [195]),
	.I2(\top/n522_48 ),
	.I3(\top/n583_15 ),
	.F(\top/n522_35 )
);
defparam \top/n522_s31 .INIT=16'h8000;
LUT4 \top/n522_s32  (
	.I0(\top/send_index [3]),
	.I1(\top/n522_81 ),
	.I2(\top/send_index [4]),
	.I3(\top/n523_117 ),
	.F(\top/n522_36 )
);
defparam \top/n522_s32 .INIT=16'h4000;
LUT4 \top/n522_s33  (
	.I0(\top/n522_61 ),
	.I1(\top/hash_out [135]),
	.I2(\top/hash_out [103]),
	.I3(\top/n522_65 ),
	.F(\top/n522_37 )
);
defparam \top/n522_s33 .INIT=16'h0777;
LUT3 \top/n522_s34  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.F(\top/n522_38 )
);
defparam \top/n522_s34 .INIT=8'h40;
LUT4 \top/n522_s35  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [95]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_52 ),
	.F(\top/n522_39 )
);
defparam \top/n522_s35 .INIT=16'h4000;
LUT3 \top/n522_s36  (
	.I0(\top/hash_out [247]),
	.I1(\top/n523_77 ),
	.I2(\top/n522_56 ),
	.F(\top/n522_40 )
);
defparam \top/n522_s36 .INIT=8'h80;
LUT4 \top/n522_s37  (
	.I0(\top/hash_out [255]),
	.I1(\top/hash_out [239]),
	.I2(\top/send_index [2]),
	.I3(\top/n522_56 ),
	.F(\top/n522_41 )
);
defparam \top/n522_s37 .INIT=16'hCA00;
LUT3 \top/n522_s38  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [139]),
	.I2(\top/n522_61 ),
	.F(\top/n522_42 )
);
defparam \top/n522_s38 .INIT=8'h80;
LUT4 \top/n522_s39  (
	.I0(\top/n522_52 ),
	.I1(\top/hash_out [75]),
	.I2(\top/hash_out [43]),
	.I3(\top/n522_45 ),
	.F(\top/n522_43 )
);
defparam \top/n522_s39 .INIT=16'h0777;
LUT2 \top/n522_s40  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [0]),
	.F(\top/n522_44 )
);
defparam \top/n522_s40 .INIT=4'h4;
LUT4 \top/n522_s41  (
	.I0(\top/send_index [3]),
	.I1(\top/send_index [6]),
	.I2(\top/send_index [5]),
	.I3(\top/send_index [4]),
	.F(\top/n522_45 )
);
defparam \top/n522_s41 .INIT=16'h1000;
LUT3 \top/n522_s42  (
	.I0(\top/hash_out [151]),
	.I1(\top/n522_61 ),
	.I2(\top/n523_77 ),
	.F(\top/n522_46 )
);
defparam \top/n522_s42 .INIT=8'h80;
LUT4 \top/n522_s43  (
	.I0(\top/hash_out [215]),
	.I1(\top/hash_out [219]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n522_47 )
);
defparam \top/n522_s43 .INIT=16'hF53F;
LUT4 \top/n522_s44  (
	.I0(\top/send_index [4]),
	.I1(\top/send_index [5]),
	.I2(\top/send_index [6]),
	.I3(\top/send_index [3]),
	.F(\top/n522_48 )
);
defparam \top/n522_s44 .INIT=16'h0100;
LUT4 \top/n522_s45  (
	.I0(\top/hash_out [171]),
	.I1(\top/send_index [1]),
	.I2(\top/n522_82 ),
	.I3(\top/n522_51 ),
	.F(\top/n522_49 )
);
defparam \top/n522_s45 .INIT=16'h2C00;
LUT4 \top/n522_s46  (
	.I0(\top/hash_out [187]),
	.I1(\top/n525_51 ),
	.I2(\top/hash_out [167]),
	.I3(\top/n522_38 ),
	.F(\top/n522_50 )
);
defparam \top/n522_s46 .INIT=16'h0777;
LUT4 \top/n522_s47  (
	.I0(\top/send_index [3]),
	.I1(\top/send_index [5]),
	.I2(\top/send_index [6]),
	.I3(\top/send_index [4]),
	.F(\top/n522_51 )
);
defparam \top/n522_s47 .INIT=16'h0100;
LUT4 \top/n522_s48  (
	.I0(\top/send_index [4]),
	.I1(\top/send_index [6]),
	.I2(\top/send_index [5]),
	.I3(\top/send_index [3]),
	.F(\top/n522_52 )
);
defparam \top/n522_s48 .INIT=16'h1000;
LUT4 \top/n522_s49  (
	.I0(\top/hash_out [67]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [1]),
	.I3(\top/n522_83 ),
	.F(\top/n522_53 )
);
defparam \top/n522_s49 .INIT=16'h00B0;
LUT4 \top/n522_s50  (
	.I0(\top/hash_out [63]),
	.I1(\top/hash_out [59]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n522_54 )
);
defparam \top/n522_s50 .INIT=16'h0C0A;
LUT4 \top/n522_s52  (
	.I0(\top/send_index [3]),
	.I1(\top/send_index [4]),
	.I2(\top/send_index [5]),
	.I3(\top/send_index [6]),
	.F(\top/n522_56 )
);
defparam \top/n522_s52 .INIT=16'h0001;
LUT3 \top/n522_s53  (
	.I0(\top/hash_out [207]),
	.I1(\top/n522_48 ),
	.I2(\top/n523_117 ),
	.F(\top/n522_57 )
);
defparam \top/n522_s53 .INIT=8'h80;
LUT4 \top/n522_s55  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [107]),
	.I2(\top/n522_65 ),
	.I3(\top/n522_44 ),
	.F(\top/n522_59 )
);
defparam \top/n522_s55 .INIT=16'h8000;
LUT4 \top/n522_s56  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [35]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_45 ),
	.F(\top/n522_60 )
);
defparam \top/n522_s56 .INIT=16'h8000;
LUT4 \top/n522_s57  (
	.I0(\top/send_index [5]),
	.I1(\top/send_index [6]),
	.I2(\top/send_index [3]),
	.I3(\top/send_index [4]),
	.F(\top/n522_61 )
);
defparam \top/n522_s57 .INIT=16'h1000;
LUT2 \top/n522_s58  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.F(\top/n522_62 )
);
defparam \top/n522_s58 .INIT=4'h1;
LUT4 \top/n522_s59  (
	.I0(\top/hash_out [111]),
	.I1(\top/send_index [0]),
	.I2(\top/n522_84 ),
	.I3(\top/send_index [2]),
	.F(\top/n522_63 )
);
defparam \top/n522_s59 .INIT=16'h2003;
LUT2 \top/n522_s60  (
	.I0(\top/n522_85 ),
	.I1(\top/send_index [0]),
	.F(\top/n522_64 )
);
defparam \top/n522_s60 .INIT=4'h4;
LUT4 \top/n522_s61  (
	.I0(\top/send_index [3]),
	.I1(\top/send_index [4]),
	.I2(\top/send_index [6]),
	.I3(\top/send_index [5]),
	.F(\top/n522_65 )
);
defparam \top/n522_s61 .INIT=16'h0100;
LUT4 \top/n522_s62  (
	.I0(\top/hash_out [231]),
	.I1(\top/send_index [1]),
	.I2(\top/n522_86 ),
	.I3(\top/n522_56 ),
	.F(\top/n522_66 )
);
defparam \top/n522_s62 .INIT=16'h8300;
LUT4 \top/n522_s63  (
	.I0(\top/hash_out [91]),
	.I1(\top/n525_51 ),
	.I2(\top/hash_out [79]),
	.I3(\top/n523_117 ),
	.F(\top/n522_67 )
);
defparam \top/n522_s63 .INIT=16'h0777;
LUT4 \top/n522_s64  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [163]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_51 ),
	.F(\top/n522_68 )
);
defparam \top/n522_s64 .INIT=16'h8000;
LUT3 \top/n522_s65  (
	.I0(\top/hash_out [199]),
	.I1(\top/n522_38 ),
	.I2(\top/n522_48 ),
	.F(\top/n522_69 )
);
defparam \top/n522_s65 .INIT=8'h80;
LUT4 \top/n522_s66  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [223]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_48 ),
	.F(\top/n522_70 )
);
defparam \top/n522_s66 .INIT=16'h4000;
LUT4 \top/n522_s67  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [143]),
	.I2(\top/n522_61 ),
	.I3(\top/n522_62 ),
	.F(\top/n522_71 )
);
defparam \top/n522_s67 .INIT=16'h8000;
LUT4 \top/n522_s68  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [191]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_51 ),
	.F(\top/n522_72 )
);
defparam \top/n522_s68 .INIT=16'h4000;
LUT4 \top/n522_s69  (
	.I0(\top/send_index [1]),
	.I1(\top/hash_out [55]),
	.I2(\top/n523_69 ),
	.I3(\top/n522_45 ),
	.F(\top/n522_73 )
);
defparam \top/n522_s69 .INIT=16'h8000;
LUT4 \top/n523_s44  (
	.I0(\top/hash_out [25]),
	.I1(\top/hash_out [17]),
	.I2(\top/send_index [0]),
	.I3(\top/n523_120 ),
	.F(\top/n523_47 )
);
defparam \top/n523_s44 .INIT=16'h5F30;
LUT4 \top/n523_s45  (
	.I0(\top/hash_out [9]),
	.I1(\top/hash_out [1]),
	.I2(\top/send_index [0]),
	.I3(\top/n523_121 ),
	.F(\top/n523_48 )
);
defparam \top/n523_s45 .INIT=16'hAFC0;
LUT4 \top/n523_s46  (
	.I0(\top/n523_122 ),
	.I1(\top/n523_123 ),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n523_49 )
);
defparam \top/n523_s46 .INIT=16'hA83F;
LUT3 \top/n523_s47  (
	.I0(\top/n523_124 ),
	.I1(\top/send_index [0]),
	.I2(\top/n522_48 ),
	.F(\top/n523_50 )
);
defparam \top/n523_s47 .INIT=8'h40;
LUT4 \top/n523_s49  (
	.I0(\top/hash_out [197]),
	.I1(\top/n522_48 ),
	.I2(\top/hash_out [69]),
	.I3(\top/n522_52 ),
	.F(\top/n523_52 )
);
defparam \top/n523_s49 .INIT=16'h0777;
LUT4 \top/n523_s50  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [189]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_51 ),
	.F(\top/n523_53 )
);
defparam \top/n523_s50 .INIT=16'h4000;
LUT3 \top/n523_s51  (
	.I0(\top/hash_out [145]),
	.I1(\top/n522_61 ),
	.I2(\top/n522_31 ),
	.F(\top/n523_54 )
);
defparam \top/n523_s51 .INIT=8'h80;
LUT4 \top/n523_s52  (
	.I0(\top/hash_out [217]),
	.I1(\top/n525_51 ),
	.I2(\top/n523_126 ),
	.I3(\top/send_index [2]),
	.F(\top/n523_55 )
);
defparam \top/n523_s52 .INIT=16'h7077;
LUT3 \top/n523_s53  (
	.I0(\top/hash_out [185]),
	.I1(\top/n522_51 ),
	.I2(\top/n525_51 ),
	.F(\top/n523_56 )
);
defparam \top/n523_s53 .INIT=8'h80;
LUT4 \top/n523_s54  (
	.I0(\top/hash_out [73]),
	.I1(\top/hash_out [65]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n523_57 )
);
defparam \top/n523_s54 .INIT=16'hCA00;
LUT3 \top/n523_s56  (
	.I0(\top/hash_out [173]),
	.I1(\top/n523_117 ),
	.I2(\top/n522_51 ),
	.F(\top/n523_59 )
);
defparam \top/n523_s56 .INIT=8'h80;
LUT4 \top/n523_s57  (
	.I0(\top/send_index [2]),
	.I1(\top/n522_62 ),
	.I2(\top/hash_out [253]),
	.I3(\top/n523_127 ),
	.F(\top/n523_60 )
);
defparam \top/n523_s57 .INIT=16'h00BF;
LUT4 \top/n523_s58  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [61]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_45 ),
	.F(\top/n523_61 )
);
defparam \top/n523_s58 .INIT=16'h4000;
LUT4 \top/n523_s59  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [129]),
	.I2(\top/n522_61 ),
	.I3(\top/n583_15 ),
	.F(\top/n523_62 )
);
defparam \top/n523_s59 .INIT=16'h8000;
LUT4 \top/n523_s60  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [225]),
	.I2(\top/n522_56 ),
	.I3(\top/n583_15 ),
	.F(\top/n523_63 )
);
defparam \top/n523_s60 .INIT=16'h8000;
LUT4 \top/n523_s61  (
	.I0(\top/send_index [1]),
	.I1(\top/hash_out [245]),
	.I2(\top/n523_128 ),
	.I3(\top/send_index [2]),
	.F(\top/n523_64 )
);
defparam \top/n523_s61 .INIT=16'hF077;
LUT4 \top/n523_s62  (
	.I0(\top/hash_out [233]),
	.I1(\top/hash_out [241]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n523_65 )
);
defparam \top/n523_s62 .INIT=16'hF53F;
LUT2 \top/n523_s63  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.F(\top/n523_66 )
);
defparam \top/n523_s63 .INIT=4'h4;
LUT4 \top/n523_s64  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [137]),
	.I2(\top/n522_61 ),
	.I3(\top/n522_44 ),
	.F(\top/n523_67 )
);
defparam \top/n523_s64 .INIT=16'h8000;
LUT4 \top/n523_s65  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [165]),
	.I2(\top/n523_66 ),
	.I3(\top/n522_51 ),
	.F(\top/n523_68 )
);
defparam \top/n523_s65 .INIT=16'h8000;
LUT2 \top/n523_s66  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [2]),
	.F(\top/n523_69 )
);
defparam \top/n523_s66 .INIT=4'h1;
LUT4 \top/n523_s67  (
	.I0(\top/hash_out [221]),
	.I1(\top/hash_out [213]),
	.I2(\top/send_index [1]),
	.I3(\top/n522_48 ),
	.F(\top/n523_70 )
);
defparam \top/n523_s67 .INIT=16'hCA00;
LUT4 \top/n523_s68  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [169]),
	.I2(\top/n522_44 ),
	.I3(\top/n522_51 ),
	.F(\top/n523_71 )
);
defparam \top/n523_s68 .INIT=16'h8000;
LUT4 \top/n523_s69  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [33]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_45 ),
	.F(\top/n523_72 )
);
defparam \top/n523_s69 .INIT=16'h8000;
LUT4 \top/n523_s70  (
	.I0(\top/n522_61 ),
	.I1(\top/hash_out [133]),
	.I2(\top/hash_out [101]),
	.I3(\top/n522_65 ),
	.F(\top/n523_73 )
);
defparam \top/n523_s70 .INIT=16'h0777;
LUT4 \top/n523_s71  (
	.I0(\top/hash_out [93]),
	.I1(\top/n522_52 ),
	.I2(\top/send_index [2]),
	.I3(\top/send_index [1]),
	.F(\top/n523_74 )
);
defparam \top/n523_s71 .INIT=16'h00F8;
LUT4 \top/n523_s72  (
	.I0(\top/hash_out [125]),
	.I1(\top/hash_out [117]),
	.I2(\top/send_index [1]),
	.I3(\top/n522_65 ),
	.F(\top/n523_75 )
);
defparam \top/n523_s72 .INIT=16'hCA00;
LUT4 \top/n523_s73  (
	.I0(\top/hash_out [177]),
	.I1(\top/hash_out [161]),
	.I2(\top/send_index [2]),
	.I3(\top/n583_15 ),
	.F(\top/n523_76 )
);
defparam \top/n523_s73 .INIT=16'hCA00;
LUT3 \top/n523_s74  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [1]),
	.F(\top/n523_77 )
);
defparam \top/n523_s74 .INIT=8'h10;
LUT4 \top/n523_s75  (
	.I0(\top/hash_out [181]),
	.I1(\top/n522_51 ),
	.I2(\top/hash_out [149]),
	.I3(\top/n522_61 ),
	.F(\top/n523_78 )
);
defparam \top/n523_s75 .INIT=16'h0777;
LUT3 \top/n523_s76  (
	.I0(\top/n523_129 ),
	.I1(\top/send_index [2]),
	.I2(\top/n522_45 ),
	.F(\top/n523_79 )
);
defparam \top/n523_s76 .INIT=8'h10;
LUT4 \top/n523_s77  (
	.I0(\top/hash_out [77]),
	.I1(\top/send_index [1]),
	.I2(\top/n523_130 ),
	.I3(\top/n522_52 ),
	.F(\top/n523_80 )
);
defparam \top/n523_s77 .INIT=16'h0E00;
LUT4 \top/n523_s78  (
	.I0(\top/hash_out [109]),
	.I1(\top/hash_out [97]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_81 )
);
defparam \top/n523_s78 .INIT=16'h3FF5;
LUT4 \top/n523_s79  (
	.I0(\top/n523_131 ),
	.I1(\top/send_index [4]),
	.I2(\top/n522_78 ),
	.I3(\top/n522_44 ),
	.F(\top/n523_82 )
);
defparam \top/n523_s79 .INIT=16'h1000;
LUT4 \top/n523_s80  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [170]),
	.I2(\top/n522_44 ),
	.I3(\top/n522_51 ),
	.F(\top/n523_83 )
);
defparam \top/n523_s80 .INIT=16'h8000;
LUT4 \top/n523_s81  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [98]),
	.I2(\top/n522_65 ),
	.I3(\top/n583_15 ),
	.F(\top/n523_84 )
);
defparam \top/n523_s81 .INIT=16'h8000;
LUT4 \top/n523_s82  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [62]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_45 ),
	.F(\top/n523_85 )
);
defparam \top/n523_s82 .INIT=16'h4000;
LUT4 \top/n523_s83  (
	.I0(\top/n522_61 ),
	.I1(\top/n523_132 ),
	.I2(\top/n523_133 ),
	.I3(\top/n522_48 ),
	.F(\top/n523_86 )
);
defparam \top/n523_s83 .INIT=16'h0777;
LUT4 \top/n523_s84  (
	.I0(\top/hash_out [158]),
	.I1(\top/hash_out [154]),
	.I2(\top/send_index [0]),
	.I3(\top/n522_61 ),
	.F(\top/n523_87 )
);
defparam \top/n523_s84 .INIT=16'hCA00;
LUT2 \top/n523_s85  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [2]),
	.F(\top/n523_88 )
);
defparam \top/n523_s85 .INIT=4'h1;
LUT4 \top/n523_s86  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [162]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_51 ),
	.F(\top/n523_89 )
);
defparam \top/n523_s86 .INIT=16'h8000;
LUT3 \top/n523_s87  (
	.I0(\top/hash_out [114]),
	.I1(\top/n522_65 ),
	.I2(\top/n522_31 ),
	.F(\top/n523_90 )
);
defparam \top/n523_s87 .INIT=8'h80;
LUT4 \top/n523_s88  (
	.I0(\top/hash_out [178]),
	.I1(\top/n522_31 ),
	.I2(\top/hash_out [174]),
	.I3(\top/n523_117 ),
	.F(\top/n523_91 )
);
defparam \top/n523_s88 .INIT=16'h0777;
LUT4 \top/n523_s89  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [106]),
	.I2(\top/n522_65 ),
	.I3(\top/n522_44 ),
	.F(\top/n523_92 )
);
defparam \top/n523_s89 .INIT=16'h8000;
LUT3 \top/n523_s90  (
	.I0(\top/hash_out [238]),
	.I1(\top/n522_56 ),
	.I2(\top/n523_117 ),
	.F(\top/n523_93 )
);
defparam \top/n523_s90 .INIT=8'h80;
LUT4 \top/n523_s91  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [234]),
	.I2(\top/n522_56 ),
	.I3(\top/n522_44 ),
	.F(\top/n523_94 )
);
defparam \top/n523_s91 .INIT=16'h8000;
LUT4 \top/n523_s92  (
	.I0(\top/hash_out [78]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/n523_134 ),
	.F(\top/n523_95 )
);
defparam \top/n523_s92 .INIT=16'hF3DF;
LUT4 \top/n523_s93  (
	.I0(\top/hash_out [94]),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [2]),
	.I3(\top/n523_135 ),
	.F(\top/n523_96 )
);
defparam \top/n523_s93 .INIT=16'h3FFD;
LUT4 \top/n523_s94  (
	.I0(\top/n522_65 ),
	.I1(\top/hash_out [122]),
	.I2(\top/hash_out [58]),
	.I3(\top/n522_45 ),
	.F(\top/n523_97 )
);
defparam \top/n523_s94 .INIT=16'h0777;
LUT4 \top/n523_s95  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [194]),
	.I2(\top/n522_48 ),
	.I3(\top/n583_15 ),
	.F(\top/n523_98 )
);
defparam \top/n523_s95 .INIT=16'h8000;
LUT4 \top/n523_s96  (
	.I0(\top/n525_51 ),
	.I1(\top/hash_out [250]),
	.I2(\top/n523_136 ),
	.I3(\top/n522_56 ),
	.F(\top/n523_99 )
);
defparam \top/n523_s96 .INIT=16'hF800;
LUT4 \top/n523_s97  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [130]),
	.I2(\top/n522_61 ),
	.I3(\top/n583_15 ),
	.F(\top/n523_100 )
);
defparam \top/n523_s97 .INIT=16'h8000;
LUT4 \top/n523_s99  (
	.I0(\top/n522_61 ),
	.I1(\top/n523_138 ),
	.I2(\top/n523_139 ),
	.I3(\top/n522_48 ),
	.F(\top/n523_102 )
);
defparam \top/n523_s99 .INIT=16'h0777;
LUT4 \top/n523_s100  (
	.I0(\top/hash_out [10]),
	.I1(\top/hash_out [2]),
	.I2(\top/send_index [0]),
	.I3(\top/n523_140 ),
	.F(\top/n523_103 )
);
defparam \top/n523_s100 .INIT=16'h305F;
LUT3 \top/n523_s101  (
	.I0(\top/hash_out [230]),
	.I1(\top/n522_38 ),
	.I2(\top/n522_56 ),
	.F(\top/n523_104 )
);
defparam \top/n523_s101 .INIT=8'h80;
LUT4 \top/n523_s102  (
	.I0(\top/hash_out [246]),
	.I1(\top/n522_56 ),
	.I2(\top/hash_out [150]),
	.I3(\top/n522_61 ),
	.F(\top/n523_105 )
);
defparam \top/n523_s102 .INIT=16'h0777;
LUT4 \top/n523_s103  (
	.I0(\top/n523_141 ),
	.I1(\top/n523_142 ),
	.I2(\top/send_index [2]),
	.I3(\top/n568_34 ),
	.F(\top/n523_106 )
);
defparam \top/n523_s103 .INIT=16'h0E00;
LUT3 \top/n523_s104  (
	.I0(\top/hash_out [110]),
	.I1(\top/n522_65 ),
	.I2(\top/n523_117 ),
	.F(\top/n523_107 )
);
defparam \top/n523_s104 .INIT=8'h80;
LUT3 \top/n523_s105  (
	.I0(\top/hash_out [186]),
	.I1(\top/n522_51 ),
	.I2(\top/n525_51 ),
	.F(\top/n523_108 )
);
defparam \top/n523_s105 .INIT=8'h80;
LUT4 \top/n523_s106  (
	.I0(\top/n525_51 ),
	.I1(\top/hash_out [218]),
	.I2(\top/n523_143 ),
	.I3(\top/n522_48 ),
	.F(\top/n523_109 )
);
defparam \top/n523_s106 .INIT=16'hF800;
LUT3 \top/n523_s107  (
	.I0(\top/n523_144 ),
	.I1(\top/send_index [0]),
	.I2(\top/n522_65 ),
	.F(\top/n523_110 )
);
defparam \top/n523_s107 .INIT=8'h10;
LUT4 \top/n523_s108  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [226]),
	.I2(\top/n522_56 ),
	.I3(\top/n583_15 ),
	.F(\top/n523_111 )
);
defparam \top/n523_s108 .INIT=16'h8000;
LUT3 \top/n523_s109  (
	.I0(\top/hash_out [146]),
	.I1(\top/n522_61 ),
	.I2(\top/n522_31 ),
	.F(\top/n523_112 )
);
defparam \top/n523_s109 .INIT=8'h80;
LUT4 \top/n523_s110  (
	.I0(\top/hash_out [38]),
	.I1(\top/hash_out [42]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_113 )
);
defparam \top/n523_s110 .INIT=16'hF53F;
LUT4 \top/n523_s111  (
	.I0(\top/hash_out [46]),
	.I1(\top/send_index [1]),
	.I2(\top/n523_145 ),
	.I3(\top/send_index [2]),
	.F(\top/n523_114 )
);
defparam \top/n523_s111 .INIT=16'hDFF3;
LUT4 \top/n523_s112  (
	.I0(\top/hash_out [206]),
	.I1(\top/hash_out [202]),
	.I2(\top/send_index [0]),
	.I3(\top/n522_48 ),
	.F(\top/n523_115 )
);
defparam \top/n523_s112 .INIT=16'hCA00;
LUT3 \top/n523_s113  (
	.I0(\top/send_index [0]),
	.I1(\top/hash_out [190]),
	.I2(\top/n522_51 ),
	.F(\top/n523_116 )
);
defparam \top/n523_s113 .INIT=8'h40;
LUT3 \top/n523_s114  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.F(\top/n523_117 )
);
defparam \top/n523_s114 .INIT=8'h10;
LUT3 \top/n523_s115  (
	.I0(\top/hash_out [90]),
	.I1(\top/n522_52 ),
	.I2(\top/n525_51 ),
	.F(\top/n523_118 )
);
defparam \top/n523_s115 .INIT=8'h80;
LUT3 \top/n523_s116  (
	.I0(\top/hash_out [210]),
	.I1(\top/n522_48 ),
	.I2(\top/n522_31 ),
	.F(\top/n523_119 )
);
defparam \top/n523_s116 .INIT=8'h80;
LUT4 \top/n525_s22  (
	.I0(\top/hash_out [184]),
	.I1(\top/hash_out [168]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n525_25 )
);
defparam \top/n525_s22 .INIT=16'h0C0A;
LUT4 \top/n525_s23  (
	.I0(\top/hash_out [172]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [0]),
	.I3(\top/n525_62 ),
	.F(\top/n525_26 )
);
defparam \top/n525_s23 .INIT=16'h0E00;
LUT4 \top/n525_s24  (
	.I0(\top/send_index [0]),
	.I1(\top/hash_out [8]),
	.I2(\top/n525_63 ),
	.I3(\top/send_index [1]),
	.F(\top/n525_27 )
);
defparam \top/n525_s24 .INIT=16'h0F77;
LUT4 \top/n525_s25  (
	.I0(\top/hash_out [20]),
	.I1(\top/hash_out [16]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n525_28 )
);
defparam \top/n525_s25 .INIT=16'hCA00;
LUT4 \top/n525_s26  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [220]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_48 ),
	.F(\top/n525_29 )
);
defparam \top/n525_s26 .INIT=16'h4000;
LUT4 \top/n525_s27  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [32]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_45 ),
	.F(\top/n525_30 )
);
defparam \top/n525_s27 .INIT=16'h8000;
LUT3 \top/n525_s28  (
	.I0(\top/n525_64 ),
	.I1(\top/send_index [1]),
	.I2(\top/n522_65 ),
	.F(\top/n525_31 )
);
defparam \top/n525_s28 .INIT=8'h10;
LUT4 \top/n525_s29  (
	.I0(\top/n522_61 ),
	.I1(\top/n525_65 ),
	.I2(\top/n525_66 ),
	.I3(\top/n568_34 ),
	.F(\top/n525_32 )
);
defparam \top/n525_s29 .INIT=16'h0777;
LUT4 \top/n525_s30  (
	.I0(\top/hash_out [128]),
	.I1(\top/send_index [0]),
	.I2(\top/n525_67 ),
	.I3(\top/send_index [2]),
	.F(\top/n525_33 )
);
defparam \top/n525_s30 .INIT=16'hB000;
LUT4 \top/n525_s31  (
	.I0(\top/n525_68 ),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [2]),
	.I3(\top/n522_65 ),
	.F(\top/n525_34 )
);
defparam \top/n525_s31 .INIT=16'h2000;
LUT4 \top/n525_s32  (
	.I0(\top/hash_out [244]),
	.I1(\top/n523_77 ),
	.I2(\top/n525_69 ),
	.I3(\top/send_index [2]),
	.F(\top/n525_35 )
);
defparam \top/n525_s32 .INIT=16'h7077;
LUT4 \top/n525_s33  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [160]),
	.I2(\top/n583_15 ),
	.I3(\top/n522_51 ),
	.F(\top/n525_36 )
);
defparam \top/n525_s33 .INIT=16'h8000;
LUT4 \top/n525_s34  (
	.I0(\top/hash_out [156]),
	.I1(\top/hash_out [136]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [2]),
	.F(\top/n525_37 )
);
defparam \top/n525_s34 .INIT=16'h3FF5;
LUT4 \top/n525_s35  (
	.I0(\top/n522_45 ),
	.I1(\top/n525_70 ),
	.I2(\top/n525_71 ),
	.I3(\top/n522_52 ),
	.F(\top/n525_38 )
);
defparam \top/n525_s35 .INIT=16'h0777;
LUT4 \top/n525_s36  (
	.I0(\top/hash_out [120]),
	.I1(\top/hash_out [96]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n525_39 )
);
defparam \top/n525_s36 .INIT=16'h3FF5;
LUT4 \top/n525_s37  (
	.I0(\top/n525_72 ),
	.I1(\top/send_index [4]),
	.I2(\top/n522_78 ),
	.I3(\top/n523_117 ),
	.F(\top/n525_40 )
);
defparam \top/n525_s37 .INIT=16'h4000;
LUT4 \top/n525_s38  (
	.I0(\top/hash_out [216]),
	.I1(\top/hash_out [200]),
	.I2(\top/send_index [2]),
	.I3(\top/n522_48 ),
	.F(\top/n525_41 )
);
defparam \top/n525_s38 .INIT=16'hCA00;
LUT3 \top/n525_s39  (
	.I0(\top/hash_out [24]),
	.I1(\top/n568_34 ),
	.I2(\top/n525_51 ),
	.F(\top/n525_42 )
);
defparam \top/n525_s39 .INIT=8'h80;
LUT4 \top/n525_s40  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [252]),
	.I2(\top/n522_56 ),
	.I3(\top/n522_62 ),
	.F(\top/n525_43 )
);
defparam \top/n525_s40 .INIT=16'h4000;
LUT4 \top/n525_s41  (
	.I0(\top/hash_out [240]),
	.I1(\top/hash_out [112]),
	.I2(\top/send_index [6]),
	.I3(\top/send_index [5]),
	.F(\top/n525_44 )
);
defparam \top/n525_s41 .INIT=16'h0C0A;
LUT4 \top/n525_s42  (
	.I0(\top/send_index [2]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [0]),
	.I3(\top/hash_out [176]),
	.F(\top/n525_45 )
);
defparam \top/n525_s42 .INIT=16'h4000;
LUT4 \top/n525_s43  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [192]),
	.I2(\top/n522_48 ),
	.I3(\top/n583_15 ),
	.F(\top/n525_46 )
);
defparam \top/n525_s43 .INIT=16'h8000;
LUT4 \top/n525_s44  (
	.I0(\top/send_index [4]),
	.I1(\top/send_index [3]),
	.I2(\top/n525_73 ),
	.I3(\top/n523_77 ),
	.F(\top/n525_47 )
);
defparam \top/n525_s44 .INIT=16'h4000;
LUT4 \top/n525_s45  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [36]),
	.I2(\top/n523_66 ),
	.I3(\top/n522_45 ),
	.F(\top/n525_48 )
);
defparam \top/n525_s45 .INIT=16'h8000;
LUT4 \top/n525_s46  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [72]),
	.I2(\top/n522_52 ),
	.I3(\top/n522_44 ),
	.F(\top/n525_49 )
);
defparam \top/n525_s46 .INIT=16'h8000;
LUT4 \top/n525_s47  (
	.I0(\top/n522_56 ),
	.I1(\top/hash_out [248]),
	.I2(\top/hash_out [56]),
	.I3(\top/n522_45 ),
	.F(\top/n525_50 )
);
defparam \top/n525_s47 .INIT=16'h0777;
LUT3 \top/n525_s48  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [0]),
	.F(\top/n525_51 )
);
defparam \top/n525_s48 .INIT=8'h10;
LUT4 \top/n525_s49  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [188]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_51 ),
	.F(\top/n525_52 )
);
defparam \top/n525_s49 .INIT=16'h4000;
LUT3 \top/n525_s50  (
	.I0(\top/hash_out [204]),
	.I1(\top/n522_48 ),
	.I2(\top/n523_117 ),
	.F(\top/n525_53 )
);
defparam \top/n525_s50 .INIT=8'h80;
LUT4 \top/n525_s51  (
	.I0(\top/hash_out [92]),
	.I1(\top/hash_out [76]),
	.I2(\top/send_index [2]),
	.I3(\top/n522_62 ),
	.F(\top/n525_54 )
);
defparam \top/n525_s51 .INIT=16'hCA00;
LUT4 \top/n525_s52  (
	.I0(\top/n583_15 ),
	.I1(\top/n525_74 ),
	.I2(\top/hash_out [88]),
	.I3(\top/n525_51 ),
	.F(\top/n525_55 )
);
defparam \top/n525_s52 .INIT=16'h0DDD;
LUT3 \top/n525_s53  (
	.I0(\top/n525_75 ),
	.I1(\top/send_index [2]),
	.I2(\top/n522_56 ),
	.F(\top/n525_56 )
);
defparam \top/n525_s53 .INIT=8'h40;
LUT4 \top/n525_s54  (
	.I0(\top/n522_61 ),
	.I1(\top/hash_out [144]),
	.I2(\top/hash_out [48]),
	.I3(\top/n522_45 ),
	.F(\top/n525_57 )
);
defparam \top/n525_s54 .INIT=16'h0777;
LUT3 \top/n525_s55  (
	.I0(\top/hash_out [196]),
	.I1(\top/n522_38 ),
	.I2(\top/n522_48 ),
	.F(\top/n525_58 )
);
defparam \top/n525_s55 .INIT=8'h80;
LUT4 \top/n525_s56  (
	.I0(\top/n522_61 ),
	.I1(\top/hash_out [148]),
	.I2(\top/hash_out [52]),
	.I3(\top/n522_45 ),
	.F(\top/n525_59 )
);
defparam \top/n525_s56 .INIT=16'h0777;
LUT4 \top/n525_s57  (
	.I0(\top/send_index [2]),
	.I1(\top/hash_out [60]),
	.I2(\top/n522_62 ),
	.I3(\top/n522_45 ),
	.F(\top/n525_60 )
);
defparam \top/n525_s57 .INIT=16'h4000;
LUT3 \top/n525_s58  (
	.I0(\top/hash_out [208]),
	.I1(\top/n522_48 ),
	.I2(\top/n522_31 ),
	.F(\top/n525_61 )
);
defparam \top/n525_s58 .INIT=8'h80;
LUT3 \top/n522_s70  (
	.I0(\top/hash_out [23]),
	.I1(\top/hash_out [19]),
	.I2(\top/send_index [0]),
	.F(\top/n522_74 )
);
defparam \top/n522_s70 .INIT=8'hCA;
LUT4 \top/n522_s71  (
	.I0(\top/hash_out [7]),
	.I1(\top/hash_out [15]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n522_75 )
);
defparam \top/n522_s71 .INIT=16'hFA0C;
LUT4 \top/n522_s72  (
	.I0(\top/hash_out [3]),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n522_76 )
);
defparam \top/n522_s72 .INIT=16'hBF00;
LUT4 \top/n522_s73  (
	.I0(\top/hash_out [115]),
	.I1(\top/hash_out [51]),
	.I2(\top/send_index [3]),
	.I3(\top/send_index [4]),
	.F(\top/n522_77 )
);
defparam \top/n522_s73 .INIT=16'h0C0A;
LUT2 \top/n522_s74  (
	.I0(\top/send_index [6]),
	.I1(\top/send_index [5]),
	.F(\top/n522_78 )
);
defparam \top/n522_s74 .INIT=4'h4;
LUT4 \top/n522_s75  (
	.I0(\top/hash_out [227]),
	.I1(\top/hash_out [131]),
	.I2(\top/send_index [3]),
	.I3(\top/send_index [4]),
	.F(\top/n522_79 )
);
defparam \top/n522_s75 .INIT=16'h3FF5;
LUT2 \top/n522_s76  (
	.I0(\top/send_index [5]),
	.I1(\top/send_index [6]),
	.F(\top/n522_80 )
);
defparam \top/n522_s76 .INIT=4'h1;
LUT4 \top/n522_s77  (
	.I0(\top/hash_out [175]),
	.I1(\top/hash_out [47]),
	.I2(\top/send_index [6]),
	.I3(\top/send_index [5]),
	.F(\top/n522_81 )
);
defparam \top/n522_s77 .INIT=16'h0C0A;
LUT4 \top/n522_s78  (
	.I0(\top/hash_out [183]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [2]),
	.F(\top/n522_82 )
);
defparam \top/n522_s78 .INIT=16'hFCC4;
LUT4 \top/n522_s79  (
	.I0(\top/hash_out [87]),
	.I1(\top/hash_out [83]),
	.I2(\top/send_index [2]),
	.I3(\top/send_index [0]),
	.F(\top/n522_83 )
);
defparam \top/n522_s79 .INIT=16'h03F5;
LUT4 \top/n522_s80  (
	.I0(\top/hash_out [127]),
	.I1(\top/hash_out [119]),
	.I2(\top/send_index [2]),
	.I3(\top/send_index [1]),
	.F(\top/n522_84 )
);
defparam \top/n522_s80 .INIT=16'h03F5;
LUT4 \top/n522_s81  (
	.I0(\top/hash_out [123]),
	.I1(\top/hash_out [99]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n522_85 )
);
defparam \top/n522_s81 .INIT=16'h3FF5;
LUT4 \top/n522_s82  (
	.I0(\top/hash_out [251]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/send_index [0]),
	.F(\top/n522_86 )
);
defparam \top/n522_s82 .INIT=16'h31F3;
LUT4 \top/n523_s117  (
	.I0(\top/hash_out [29]),
	.I1(\top/hash_out [21]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_120 )
);
defparam \top/n523_s117 .INIT=16'h03F5;
LUT4 \top/n523_s118  (
	.I0(\top/hash_out [13]),
	.I1(\top/hash_out [5]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_121 )
);
defparam \top/n523_s118 .INIT=16'h0CFA;
LUT4 \top/n523_s119  (
	.I0(\top/hash_out [37]),
	.I1(\top/hash_out [41]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_122 )
);
defparam \top/n523_s119 .INIT=16'hF53F;
LUT4 \top/n523_s120  (
	.I0(\top/hash_out [45]),
	.I1(\top/hash_out [49]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n523_123 )
);
defparam \top/n523_s120 .INIT=16'hCF05;
LUT4 \top/n523_s121  (
	.I0(\top/hash_out [201]),
	.I1(\top/hash_out [209]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n523_124 )
);
defparam \top/n523_s121 .INIT=16'hF53F;
LUT3 \top/n523_s122  (
	.I0(\top/hash_out [157]),
	.I1(\top/hash_out [141]),
	.I2(\top/send_index [2]),
	.F(\top/n523_125 )
);
defparam \top/n523_s122 .INIT=8'h35;
LUT4 \top/n523_s123  (
	.I0(\top/hash_out [205]),
	.I1(\top/hash_out [193]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_126 )
);
defparam \top/n523_s123 .INIT=16'h3FF5;
LUT4 \top/n523_s124  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [0]),
	.I3(\top/hash_out [249]),
	.F(\top/n523_127 )
);
defparam \top/n523_s124 .INIT=16'h1000;
LUT3 \top/n523_s125  (
	.I0(\top/hash_out [237]),
	.I1(\top/hash_out [229]),
	.I2(\top/send_index [1]),
	.F(\top/n523_128 )
);
defparam \top/n523_s125 .INIT=8'h35;
LUT4 \top/n523_s126  (
	.I0(\top/hash_out [53]),
	.I1(\top/hash_out [57]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_129 )
);
defparam \top/n523_s126 .INIT=16'hF53F;
LUT4 \top/n523_s127  (
	.I0(\top/hash_out [81]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_130 )
);
defparam \top/n523_s127 .INIT=16'hDFF3;
LUT4 \top/n523_s128  (
	.I0(\top/hash_out [89]),
	.I1(\top/hash_out [105]),
	.I2(\top/send_index [2]),
	.I3(\top/send_index [3]),
	.F(\top/n523_131 )
);
defparam \top/n523_s128 .INIT=16'hF53F;
LUT4 \top/n523_s129  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [134]),
	.F(\top/n523_132 )
);
defparam \top/n523_s129 .INIT=16'h4000;
LUT4 \top/n523_s130  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [1]),
	.I3(\top/hash_out [214]),
	.F(\top/n523_133 )
);
defparam \top/n523_s130 .INIT=16'h1000;
LUT4 \top/n523_s131  (
	.I0(\top/hash_out [82]),
	.I1(\top/hash_out [86]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n523_134 )
);
defparam \top/n523_s131 .INIT=16'hAFC0;
LUT4 \top/n523_s132  (
	.I0(\top/hash_out [66]),
	.I1(\top/hash_out [74]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_135 )
);
defparam \top/n523_s132 .INIT=16'hAFC0;
LUT4 \top/n523_s133  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [254]),
	.F(\top/n523_136 )
);
defparam \top/n523_s133 .INIT=16'h0100;
LUT3 \top/n523_s134  (
	.I0(\top/hash_out [182]),
	.I1(\top/hash_out [166]),
	.I2(\top/send_index [2]),
	.F(\top/n523_137 )
);
defparam \top/n523_s134 .INIT=8'hCA;
LUT4 \top/n523_s135  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [138]),
	.F(\top/n523_138 )
);
defparam \top/n523_s135 .INIT=16'h4000;
LUT4 \top/n523_s136  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [222]),
	.F(\top/n523_139 )
);
defparam \top/n523_s136 .INIT=16'h0100;
LUT4 \top/n523_s137  (
	.I0(\top/hash_out [6]),
	.I1(\top/hash_out [14]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_140 )
);
defparam \top/n523_s137 .INIT=16'hFA0C;
LUT4 \top/n523_s138  (
	.I0(\top/hash_out [30]),
	.I1(\top/hash_out [26]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n523_141 )
);
defparam \top/n523_s138 .INIT=16'h0C0A;
LUT4 \top/n523_s139  (
	.I0(\top/hash_out [22]),
	.I1(\top/hash_out [18]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_142 )
);
defparam \top/n523_s139 .INIT=16'hCA00;
LUT4 \top/n523_s140  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [198]),
	.F(\top/n523_143 )
);
defparam \top/n523_s140 .INIT=16'h4000;
LUT4 \top/n523_s141  (
	.I0(\top/hash_out [126]),
	.I1(\top/hash_out [102]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n523_144 )
);
defparam \top/n523_s141 .INIT=16'h3FF5;
LUT4 \top/n523_s142  (
	.I0(\top/hash_out [54]),
	.I1(\top/hash_out [50]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n523_145 )
);
defparam \top/n523_s142 .INIT=16'h305F;
LUT4 \top/n525_s59  (
	.I0(\top/hash_out [164]),
	.I1(\top/hash_out [180]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [2]),
	.F(\top/n525_62 )
);
defparam \top/n525_s59 .INIT=16'hAFC0;
LUT3 \top/n525_s60  (
	.I0(\top/hash_out [4]),
	.I1(\top/hash_out [0]),
	.I2(\top/send_index [0]),
	.F(\top/n525_63 )
);
defparam \top/n525_s60 .INIT=8'hCA;
LUT4 \top/n525_s61  (
	.I0(\top/hash_out [124]),
	.I1(\top/hash_out [104]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [2]),
	.F(\top/n525_64 )
);
defparam \top/n525_s61 .INIT=16'h3FF5;
LUT4 \top/n525_s62  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [0]),
	.I3(\top/hash_out [152]),
	.F(\top/n525_65 )
);
defparam \top/n525_s62 .INIT=16'h1000;
LUT4 \top/n525_s63  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [28]),
	.F(\top/n525_66 )
);
defparam \top/n525_s63 .INIT=16'h0100;
LUT4 \top/n525_s64  (
	.I0(\top/hash_out [132]),
	.I1(\top/hash_out [140]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n525_67 )
);
defparam \top/n525_s64 .INIT=16'hFA0C;
LUT3 \top/n525_s65  (
	.I0(\top/hash_out [108]),
	.I1(\top/hash_out [100]),
	.I2(\top/send_index [1]),
	.F(\top/n525_68 )
);
defparam \top/n525_s65 .INIT=8'hCA;
LUT4 \top/n525_s66  (
	.I0(\top/hash_out [236]),
	.I1(\top/hash_out [224]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n525_69 )
);
defparam \top/n525_s66 .INIT=16'h3FF5;
LUT4 \top/n525_s67  (
	.I0(\top/send_index [1]),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [40]),
	.F(\top/n525_70 )
);
defparam \top/n525_s67 .INIT=16'h4000;
LUT4 \top/n525_s68  (
	.I0(\top/send_index [0]),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/hash_out [68]),
	.F(\top/n525_71 )
);
defparam \top/n525_s68 .INIT=16'h4000;
LUT3 \top/n525_s69  (
	.I0(\top/hash_out [44]),
	.I1(\top/hash_out [12]),
	.I2(\top/send_index [3]),
	.F(\top/n525_72 )
);
defparam \top/n525_s69 .INIT=8'h35;
LUT4 \top/n525_s70  (
	.I0(\top/hash_out [212]),
	.I1(\top/hash_out [84]),
	.I2(\top/send_index [6]),
	.I3(\top/send_index [5]),
	.F(\top/n525_73 )
);
defparam \top/n525_s70 .INIT=16'h0C0A;
LUT3 \top/n525_s71  (
	.I0(\top/hash_out [80]),
	.I1(\top/hash_out [64]),
	.I2(\top/send_index [2]),
	.F(\top/n525_74 )
);
defparam \top/n525_s71 .INIT=8'h35;
LUT4 \top/n525_s72  (
	.I0(\top/hash_out [228]),
	.I1(\top/hash_out [232]),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n525_75 )
);
defparam \top/n525_s72 .INIT=16'hF53F;
LUT4 \top/n524_s1  (
	.I0(\top/n523_6 ),
	.I1(\top/n523_5 ),
	.I2(\top/n522_5 ),
	.I3(\top/n525_4 ),
	.F(\top/n524_5 )
);
defparam \top/n524_s1 .INIT=16'h3433;
LUT4 \top/n523_s143  (
	.I0(\top/n522_5 ),
	.I1(\top/n525_4 ),
	.I2(\top/n523_5 ),
	.I3(\top/n523_6 ),
	.F(\top/n523_147 )
);
defparam \top/n523_s143 .INIT=16'h00BF;
LUT4 \top/n570_s6  (
	.I0(\top/tx_busy_Z ),
	.I1(\top/state [2]),
	.I2(\top/state [1]),
	.I3(\top/state [0]),
	.F(\top/n570_11 )
);
defparam \top/n570_s6 .INIT=16'h1000;
LUT4 \top/tx_data_4_s10  (
	.I0(\top/n522_5 ),
	.I1(\top/n525_4 ),
	.I2(\top/tx_data_4_15 ),
	.I3(\top/n636_5 ),
	.F(\top/tx_data_4_19 )
);
defparam \top/tx_data_4_s10 .INIT=16'h00FE;
LUT4 \top/tx_data_5_s11  (
	.I0(\top/n636_5 ),
	.I1(\top/tx_data_4_15 ),
	.I2(\top/n522_5 ),
	.I3(\top/n525_4 ),
	.F(\top/tx_data_5_19 )
);
defparam \top/tx_data_5_s11 .INIT=16'hEEEF;
LUT3 \top/n603_s4  (
	.I0(\top/state [1]),
	.I1(\top/state [2]),
	.I2(\top/n568_26 ),
	.F(\top/n603_10 )
);
defparam \top/n603_s4 .INIT=8'h10;
LUT4 \top/n586_s7  (
	.I0(\top/rx_valid_Z ),
	.I1(\top/state [0]),
	.I2(\top/state [1]),
	.I3(\top/state [2]),
	.F(\top/n586_12 )
);
defparam \top/n586_s7 .INIT=16'h0008;
LUT4 \top/n523_s144  (
	.I0(\top/n523_137 ),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [1]),
	.I3(\top/n522_51 ),
	.F(\top/n523_149 )
);
defparam \top/n523_s144 .INIT=16'h2000;
LUT4 \top/n525_s73  (
	.I0(\top/n523_6 ),
	.I1(\top/n523_5 ),
	.I2(\top/n522_5 ),
	.I3(\top/n525_4 ),
	.F(\top/n525_77 )
);
defparam \top/n525_s73 .INIT=16'h07F8;
LUT4 \top/n522_s84  (
	.I0(\top/n522_61 ),
	.I1(\top/send_index [1]),
	.I2(\top/send_index [2]),
	.I3(\top/send_index [0]),
	.F(\top/n522_90 )
);
defparam \top/n522_s84 .INIT=16'h0200;
LUT4 \top/n523_s145  (
	.I0(\top/hash_out [121]),
	.I1(\top/n522_65 ),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n523_151 )
);
defparam \top/n523_s145 .INIT=16'h0800;
LUT4 \top/n522_s85  (
	.I0(\top/hash_out [203]),
	.I1(\top/n522_48 ),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n522_92 )
);
defparam \top/n522_s85 .INIT=16'h0800;
LUT4 \top/n522_s86  (
	.I0(\top/n522_43 ),
	.I1(\top/send_index [2]),
	.I2(\top/send_index [1]),
	.I3(\top/send_index [0]),
	.F(\top/n522_94 )
);
defparam \top/n522_s86 .INIT=16'h0400;
LUT4 \top/n523_s146  (
	.I0(\top/n523_125 ),
	.I1(\top/n522_61 ),
	.I2(\top/send_index [0]),
	.I3(\top/send_index [1]),
	.F(\top/n523_153 )
);
defparam \top/n523_s146 .INIT=16'h0004;
LUT3 \top/n582_s11  (
	.I0(\top/send_index [2]),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [1]),
	.F(\top/n582_17 )
);
defparam \top/n582_s11 .INIT=8'h80;
LUT4 \top/n583_s11  (
	.I0(\top/send_index [2]),
	.I1(\top/send_index [0]),
	.I2(\top/send_index [1]),
	.I3(\top/state [0]),
	.F(\top/n583_17 )
);
defparam \top/n583_s11 .INIT=16'h6A00;
LUT4 \top/n569_s16  (
	.I0(\top/state [0]),
	.I1(\top/state [2]),
	.I2(\top/state_0_9 ),
	.I3(\top/n568_25 ),
	.F(\top/n569_27 )
);
defparam \top/n569_s16 .INIT=16'h19AA;
LUT3 \top/state_0_s6  (
	.I0(\top/state [2]),
	.I1(\top/state_0_9 ),
	.I2(\top/n568_25 ),
	.F(\top/state_0_13 )
);
defparam \top/state_0_s6 .INIT=8'hD0;
LUT3 \top/n522_s87  (
	.I0(\top/n522_5 ),
	.I1(\top/n523_6 ),
	.I2(\top/n523_5 ),
	.F(\top/n522_96 )
);
defparam \top/n522_s87 .INIT=8'h40;
DFFC \top/data_valid_s0  (
	.D(\top/n586_12 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/data_valid )
);
defparam \top/data_valid_s0 .INIT=1'b0;
DFFC \top/data_last_s0  (
	.D(\top/n603_10 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/data_last )
);
defparam \top/data_last_s0 .INIT=1'b0;
DFFC \top/tx_start_s0  (
	.D(\top/n570_11 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/tx_start )
);
defparam \top/tx_start_s0 .INIT=1'b0;
DFFCE \top/send_index_6_s0  (
	.D(\top/n579_15 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [6])
);
defparam \top/send_index_6_s0 .INIT=1'b0;
DFFCE \top/send_index_5_s0  (
	.D(\top/n580_14 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [5])
);
defparam \top/send_index_5_s0 .INIT=1'b0;
DFFCE \top/send_index_4_s0  (
	.D(\top/n581_14 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [4])
);
defparam \top/send_index_4_s0 .INIT=1'b0;
DFFCE \top/send_index_3_s0  (
	.D(\top/n582_14 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [3])
);
defparam \top/send_index_3_s0 .INIT=1'b0;
DFFCE \top/send_index_2_s0  (
	.D(\top/n583_17 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [2])
);
defparam \top/send_index_2_s0 .INIT=1'b0;
DFFCE \top/send_index_1_s0  (
	.D(\top/n584_14 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [1])
);
defparam \top/send_index_1_s0 .INIT=1'b0;
DFFCE \top/send_index_0_s0  (
	.D(\top/n585_15 ),
	.CLK(clk),
	.CE(\top/send_index_6_7 ),
	.CLEAR(rst),
	.Q(\top/send_index [0])
);
defparam \top/send_index_0_s0 .INIT=1'b0;
DFFE \top/tx_data_6_s0  (
	.D(\top/n636_5 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [6])
);
defparam \top/tx_data_6_s0 .INIT=1'b0;
DFFE \top/tx_data_3_s0  (
	.D(\top/n522_96 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [3])
);
defparam \top/tx_data_3_s0 .INIT=1'b0;
DFFE \top/tx_data_2_s0  (
	.D(\top/n523_147 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [2])
);
defparam \top/tx_data_2_s0 .INIT=1'b0;
DFFE \top/tx_data_1_s0  (
	.D(\top/n524_5 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [1])
);
defparam \top/tx_data_1_s0 .INIT=1'b0;
DFFE \top/tx_data_0_s0  (
	.D(\top/n525_77 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [0])
);
defparam \top/tx_data_0_s0 .INIT=1'b0;
DFFE \top/data_in_7_s0  (
	.D(\top/rx_data_Z [7]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [7])
);
defparam \top/data_in_7_s0 .INIT=1'b0;
DFFE \top/data_in_6_s0  (
	.D(\top/rx_data_Z [6]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [6])
);
defparam \top/data_in_6_s0 .INIT=1'b0;
DFFE \top/data_in_5_s0  (
	.D(\top/rx_data_Z [5]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [5])
);
defparam \top/data_in_5_s0 .INIT=1'b0;
DFFE \top/data_in_4_s0  (
	.D(\top/rx_data_Z [4]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [4])
);
defparam \top/data_in_4_s0 .INIT=1'b0;
DFFE \top/data_in_3_s0  (
	.D(\top/rx_data_Z [3]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [3])
);
defparam \top/data_in_3_s0 .INIT=1'b0;
DFFE \top/data_in_2_s0  (
	.D(\top/rx_data_Z [2]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [2])
);
defparam \top/data_in_2_s0 .INIT=1'b0;
DFFE \top/data_in_1_s0  (
	.D(\top/rx_data_Z [1]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [1])
);
defparam \top/data_in_1_s0 .INIT=1'b0;
DFFE \top/data_in_0_s0  (
	.D(\top/rx_data_Z [0]),
	.CLK(clk),
	.CE(\top/data_in_7_6 ),
	.Q(\top/data_in [0])
);
defparam \top/data_in_0_s0 .INIT=1'b0;
DFFCE \top/state_2_s1  (
	.D(\top/n567_20 ),
	.CLK(clk),
	.CE(\top/state_0_13 ),
	.CLEAR(rst),
	.Q(\top/state [2])
);
defparam \top/state_2_s1 .INIT=1'b0;
DFFE \top/tx_data_4_s6  (
	.D(\top/tx_data_4_19 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [4])
);
defparam \top/tx_data_4_s6 .INIT=1'b0;
DFFE \top/tx_data_5_s6  (
	.D(\top/tx_data_5_19 ),
	.CLK(clk),
	.CE(\top/tx_data_4_15 ),
	.Q(\top/tx_data [5])
);
defparam \top/tx_data_5_s6 .INIT=1'b0;
DFFCE \top/state_1_s1  (
	.D(\top/n568_23 ),
	.CLK(clk),
	.CE(\top/n568_25 ),
	.CLEAR(rst),
	.Q(\top/state [1])
);
defparam \top/state_1_s1 .INIT=1'b0;
DFFC \top/state_0_s5  (
	.D(\top/n569_27 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/state [0])
);
defparam \top/state_0_s5 .INIT=1'b0;
LUT2 \top/uart_rx_inst/n200_s6  (
	.I0(\top/uart_rx_inst/state [0]),
	.I1(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n200_12 )
);
defparam \top/uart_rx_inst/n200_s6 .INIT=4'h6;
LUT3 \top/uart_rx_inst/n191_s5  (
	.I0(\top/uart_rx_inst/state [0]),
	.I1(\top/uart_rx_inst/state [1]),
	.I2(\top/uart_rx_inst/n191_10 ),
	.F(\top/uart_rx_inst/n191_9 )
);
defparam \top/uart_rx_inst/n191_s5 .INIT=8'h80;
LUT4 \top/uart_rx_inst/bit_cnt_3_s3  (
	.I0(\top/uart_rx_inst/n191_10 ),
	.I1(\top/uart_rx_inst/rx_dd ),
	.I2(\top/uart_rx_inst/state [0]),
	.I3(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/bit_cnt_3_8 )
);
defparam \top/uart_rx_inst/bit_cnt_3_s3 .INIT=16'h0A03;
LUT4 \top/uart_rx_inst/state_0_s4  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/rx_dd ),
	.I2(\top/uart_rx_inst/n191_10 ),
	.I3(\top/uart_rx_inst/state_0_10 ),
	.F(\top/uart_rx_inst/n139_4 )
);
defparam \top/uart_rx_inst/state_0_s4 .INIT=16'h11F0;
LUT2 \top/uart_rx_inst/n217_s6  (
	.I0(\top/uart_rx_inst/baud_cnt [0]),
	.I1(\top/uart_rx_inst/n217_14 ),
	.F(\top/uart_rx_inst/n217_11 )
);
defparam \top/uart_rx_inst/n217_s6 .INIT=4'h4;
LUT4 \top/uart_rx_inst/n215_s6  (
	.I0(\top/uart_rx_inst/baud_cnt [0]),
	.I1(\top/uart_rx_inst/baud_cnt [1]),
	.I2(\top/uart_rx_inst/n217_14 ),
	.I3(\top/uart_rx_inst/baud_cnt [2]),
	.F(\top/uart_rx_inst/n215_11 )
);
defparam \top/uart_rx_inst/n215_s6 .INIT=16'h7080;
LUT3 \top/uart_rx_inst/n214_s6  (
	.I0(\top/uart_rx_inst/n217_14 ),
	.I1(\top/uart_rx_inst/baud_cnt [3]),
	.I2(\top/uart_rx_inst/n214_12 ),
	.F(\top/uart_rx_inst/n214_11 )
);
defparam \top/uart_rx_inst/n214_s6 .INIT=8'h28;
LUT3 \top/uart_rx_inst/n211_s6  (
	.I0(\top/uart_rx_inst/n217_14 ),
	.I1(\top/uart_rx_inst/baud_cnt [6]),
	.I2(\top/uart_rx_inst/n211_12 ),
	.F(\top/uart_rx_inst/n211_11 )
);
defparam \top/uart_rx_inst/n211_s6 .INIT=8'h28;
LUT3 \top/uart_rx_inst/n208_s6  (
	.I0(\top/uart_rx_inst/n217_14 ),
	.I1(\top/uart_rx_inst/baud_cnt [9]),
	.I2(\top/uart_rx_inst/n208_12 ),
	.F(\top/uart_rx_inst/n208_11 )
);
defparam \top/uart_rx_inst/n208_s6 .INIT=8'h28;
LUT4 \top/uart_rx_inst/n207_s6  (
	.I0(\top/uart_rx_inst/baud_cnt [9]),
	.I1(\top/uart_rx_inst/n208_12 ),
	.I2(\top/uart_rx_inst/n217_14 ),
	.I3(\top/uart_rx_inst/baud_cnt [10]),
	.F(\top/uart_rx_inst/n207_11 )
);
defparam \top/uart_rx_inst/n207_s6 .INIT=16'h7080;
LUT3 \top/uart_rx_inst/n206_s6  (
	.I0(\top/uart_rx_inst/n217_14 ),
	.I1(\top/uart_rx_inst/baud_cnt [11]),
	.I2(\top/uart_rx_inst/n206_12 ),
	.F(\top/uart_rx_inst/n206_11 )
);
defparam \top/uart_rx_inst/n206_s6 .INIT=8'h28;
LUT4 \top/uart_rx_inst/n205_s6  (
	.I0(\top/uart_rx_inst/baud_cnt [11]),
	.I1(\top/uart_rx_inst/n206_12 ),
	.I2(\top/uart_rx_inst/n217_14 ),
	.I3(\top/uart_rx_inst/baud_cnt [12]),
	.F(\top/uart_rx_inst/n205_11 )
);
defparam \top/uart_rx_inst/n205_s6 .INIT=16'h7080;
LUT3 \top/uart_rx_inst/n204_s6  (
	.I0(\top/uart_rx_inst/n217_14 ),
	.I1(\top/uart_rx_inst/n204_12 ),
	.I2(\top/uart_rx_inst/baud_cnt [13]),
	.F(\top/uart_rx_inst/n204_11 )
);
defparam \top/uart_rx_inst/n204_s6 .INIT=8'h28;
LUT3 \top/uart_rx_inst/n203_s6  (
	.I0(\top/uart_rx_inst/n217_14 ),
	.I1(\top/uart_rx_inst/baud_cnt [14]),
	.I2(\top/uart_rx_inst/n203_12 ),
	.F(\top/uart_rx_inst/n203_11 )
);
defparam \top/uart_rx_inst/n203_s6 .INIT=8'h28;
LUT4 \top/uart_rx_inst/n202_s6  (
	.I0(\top/uart_rx_inst/baud_cnt [14]),
	.I1(\top/uart_rx_inst/n203_12 ),
	.I2(\top/uart_rx_inst/n217_14 ),
	.I3(\top/uart_rx_inst/baud_cnt [15]),
	.F(\top/uart_rx_inst/n202_11 )
);
defparam \top/uart_rx_inst/n202_s6 .INIT=16'h7080;
LUT2 \top/uart_rx_inst/n229_s7  (
	.I0(\top/uart_rx_inst/bit_cnt [0]),
	.I1(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n229_12 )
);
defparam \top/uart_rx_inst/n229_s7 .INIT=4'h4;
LUT3 \top/uart_rx_inst/n228_s6  (
	.I0(\top/uart_rx_inst/bit_cnt [0]),
	.I1(\top/uart_rx_inst/bit_cnt [1]),
	.I2(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n228_11 )
);
defparam \top/uart_rx_inst/n228_s6 .INIT=8'h60;
LUT4 \top/uart_rx_inst/n227_s6  (
	.I0(\top/uart_rx_inst/bit_cnt [0]),
	.I1(\top/uart_rx_inst/bit_cnt [1]),
	.I2(\top/uart_rx_inst/bit_cnt [2]),
	.I3(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n227_11 )
);
defparam \top/uart_rx_inst/n227_s6 .INIT=16'h7800;
LUT3 \top/uart_rx_inst/n226_s6  (
	.I0(\top/uart_rx_inst/n226_12 ),
	.I1(\top/uart_rx_inst/bit_cnt [3]),
	.I2(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n226_11 )
);
defparam \top/uart_rx_inst/n226_s6 .INIT=8'h60;
LUT2 \top/uart_rx_inst/n225_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [1]),
	.F(\top/uart_rx_inst/n225_11 )
);
defparam \top/uart_rx_inst/n225_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n224_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [2]),
	.F(\top/uart_rx_inst/n224_11 )
);
defparam \top/uart_rx_inst/n224_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n223_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [3]),
	.F(\top/uart_rx_inst/n223_11 )
);
defparam \top/uart_rx_inst/n223_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n222_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [4]),
	.F(\top/uart_rx_inst/n222_11 )
);
defparam \top/uart_rx_inst/n222_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n221_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [5]),
	.F(\top/uart_rx_inst/n221_11 )
);
defparam \top/uart_rx_inst/n221_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n220_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [6]),
	.F(\top/uart_rx_inst/n220_11 )
);
defparam \top/uart_rx_inst/n220_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n219_s6  (
	.I0(\top/uart_rx_inst/state [1]),
	.I1(\top/uart_rx_inst/shift_reg [7]),
	.F(\top/uart_rx_inst/n219_11 )
);
defparam \top/uart_rx_inst/n219_s6 .INIT=4'h8;
LUT2 \top/uart_rx_inst/n218_s7  (
	.I0(\top/uart_rx_inst/rx_dd ),
	.I1(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n218_12 )
);
defparam \top/uart_rx_inst/n218_s7 .INIT=4'h8;
LUT4 \top/uart_rx_inst/n19_s2  (
	.I0(\top/uart_rx_inst/baud_cnt [3]),
	.I1(\top/uart_rx_inst/n214_12 ),
	.I2(\top/uart_rx_inst/baud_cnt_15_9 ),
	.I3(\top/uart_rx_inst/baud_cnt [4]),
	.F(\top/uart_rx_inst/n19_6 )
);
defparam \top/uart_rx_inst/n19_s2 .INIT=16'hF7F8;
LUT4 \top/uart_rx_inst/n18_s2  (
	.I0(\top/uart_rx_inst/baud_cnt_15_9 ),
	.I1(\top/uart_rx_inst/n191_10 ),
	.I2(\top/uart_rx_inst/n18_7 ),
	.I3(\top/uart_rx_inst/baud_cnt [5]),
	.F(\top/uart_rx_inst/n18_6 )
);
defparam \top/uart_rx_inst/n18_s2 .INIT=16'hABBA;
LUT4 \top/uart_rx_inst/n16_s2  (
	.I0(\top/uart_rx_inst/baud_cnt [6]),
	.I1(\top/uart_rx_inst/n211_12 ),
	.I2(\top/uart_rx_inst/baud_cnt_15_9 ),
	.I3(\top/uart_rx_inst/baud_cnt [7]),
	.F(\top/uart_rx_inst/n16_6 )
);
defparam \top/uart_rx_inst/n16_s2 .INIT=16'hF7F8;
LUT4 \top/uart_rx_inst/n15_s2  (
	.I0(\top/uart_rx_inst/baud_cnt_15_9 ),
	.I1(\top/uart_rx_inst/n191_10 ),
	.I2(\top/uart_rx_inst/n15_7 ),
	.I3(\top/uart_rx_inst/baud_cnt [8]),
	.F(\top/uart_rx_inst/n15_6 )
);
defparam \top/uart_rx_inst/n15_s2 .INIT=16'hABBA;
LUT4 \top/uart_rx_inst/n191_s6  (
	.I0(\top/uart_rx_inst/n191_11 ),
	.I1(\top/uart_rx_inst/n191_12 ),
	.I2(\top/uart_rx_inst/n191_13 ),
	.I3(\top/uart_rx_inst/n191_14 ),
	.F(\top/uart_rx_inst/n191_10 )
);
defparam \top/uart_rx_inst/n191_s6 .INIT=16'h8000;
LUT2 \top/uart_rx_inst/baud_cnt_15_s4  (
	.I0(\top/uart_rx_inst/state [0]),
	.I1(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/baud_cnt_15_9 )
);
defparam \top/uart_rx_inst/baud_cnt_15_s4 .INIT=4'h1;
LUT3 \top/uart_rx_inst/state_0_s5  (
	.I0(\top/uart_rx_inst/state_0_11 ),
	.I1(\top/uart_rx_inst/state [1]),
	.I2(\top/uart_rx_inst/state [0]),
	.F(\top/uart_rx_inst/state_0_10 )
);
defparam \top/uart_rx_inst/state_0_s5 .INIT=8'h07;
LUT3 \top/uart_rx_inst/n214_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [0]),
	.I1(\top/uart_rx_inst/baud_cnt [1]),
	.I2(\top/uart_rx_inst/baud_cnt [2]),
	.F(\top/uart_rx_inst/n214_12 )
);
defparam \top/uart_rx_inst/n214_s7 .INIT=8'h80;
LUT4 \top/uart_rx_inst/n211_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [3]),
	.I1(\top/uart_rx_inst/baud_cnt [4]),
	.I2(\top/uart_rx_inst/baud_cnt [5]),
	.I3(\top/uart_rx_inst/n214_12 ),
	.F(\top/uart_rx_inst/n211_12 )
);
defparam \top/uart_rx_inst/n211_s7 .INIT=16'h8000;
LUT4 \top/uart_rx_inst/n208_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [6]),
	.I1(\top/uart_rx_inst/baud_cnt [7]),
	.I2(\top/uart_rx_inst/baud_cnt [8]),
	.I3(\top/uart_rx_inst/n211_12 ),
	.F(\top/uart_rx_inst/n208_12 )
);
defparam \top/uart_rx_inst/n208_s7 .INIT=16'h8000;
LUT3 \top/uart_rx_inst/n206_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [9]),
	.I1(\top/uart_rx_inst/baud_cnt [10]),
	.I2(\top/uart_rx_inst/n208_12 ),
	.F(\top/uart_rx_inst/n206_12 )
);
defparam \top/uart_rx_inst/n206_s7 .INIT=8'h80;
LUT3 \top/uart_rx_inst/n204_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [11]),
	.I1(\top/uart_rx_inst/baud_cnt [12]),
	.I2(\top/uart_rx_inst/n206_12 ),
	.F(\top/uart_rx_inst/n204_12 )
);
defparam \top/uart_rx_inst/n204_s7 .INIT=8'h80;
LUT4 \top/uart_rx_inst/n203_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [11]),
	.I1(\top/uart_rx_inst/baud_cnt [12]),
	.I2(\top/uart_rx_inst/baud_cnt [13]),
	.I3(\top/uart_rx_inst/n206_12 ),
	.F(\top/uart_rx_inst/n203_12 )
);
defparam \top/uart_rx_inst/n203_s7 .INIT=16'h8000;
LUT3 \top/uart_rx_inst/n226_s7  (
	.I0(\top/uart_rx_inst/bit_cnt [0]),
	.I1(\top/uart_rx_inst/bit_cnt [1]),
	.I2(\top/uart_rx_inst/bit_cnt [2]),
	.F(\top/uart_rx_inst/n226_12 )
);
defparam \top/uart_rx_inst/n226_s7 .INIT=8'h80;
LUT3 \top/uart_rx_inst/n18_s3  (
	.I0(\top/uart_rx_inst/baud_cnt [3]),
	.I1(\top/uart_rx_inst/baud_cnt [4]),
	.I2(\top/uart_rx_inst/n214_12 ),
	.F(\top/uart_rx_inst/n18_7 )
);
defparam \top/uart_rx_inst/n18_s3 .INIT=8'h80;
LUT3 \top/uart_rx_inst/n15_s3  (
	.I0(\top/uart_rx_inst/baud_cnt [6]),
	.I1(\top/uart_rx_inst/baud_cnt [7]),
	.I2(\top/uart_rx_inst/n211_12 ),
	.F(\top/uart_rx_inst/n15_7 )
);
defparam \top/uart_rx_inst/n15_s3 .INIT=8'h80;
LUT4 \top/uart_rx_inst/n191_s7  (
	.I0(\top/uart_rx_inst/baud_cnt [10]),
	.I1(\top/uart_rx_inst/baud_cnt [11]),
	.I2(\top/uart_rx_inst/baud_cnt [8]),
	.I3(\top/uart_rx_inst/baud_cnt [9]),
	.F(\top/uart_rx_inst/n191_11 )
);
defparam \top/uart_rx_inst/n191_s7 .INIT=16'h1000;
LUT4 \top/uart_rx_inst/n191_s8  (
	.I0(\top/uart_rx_inst/baud_cnt [0]),
	.I1(\top/uart_rx_inst/baud_cnt [1]),
	.I2(\top/uart_rx_inst/baud_cnt [5]),
	.I3(\top/uart_rx_inst/baud_cnt [6]),
	.F(\top/uart_rx_inst/n191_12 )
);
defparam \top/uart_rx_inst/n191_s8 .INIT=16'h1000;
LUT4 \top/uart_rx_inst/n191_s9  (
	.I0(\top/uart_rx_inst/baud_cnt [12]),
	.I1(\top/uart_rx_inst/baud_cnt [13]),
	.I2(\top/uart_rx_inst/baud_cnt [14]),
	.I3(\top/uart_rx_inst/baud_cnt [15]),
	.F(\top/uart_rx_inst/n191_13 )
);
defparam \top/uart_rx_inst/n191_s9 .INIT=16'h0001;
LUT4 \top/uart_rx_inst/n191_s10  (
	.I0(\top/uart_rx_inst/baud_cnt [3]),
	.I1(\top/uart_rx_inst/baud_cnt [4]),
	.I2(\top/uart_rx_inst/baud_cnt [7]),
	.I3(\top/uart_rx_inst/baud_cnt [2]),
	.F(\top/uart_rx_inst/n191_14 )
);
defparam \top/uart_rx_inst/n191_s10 .INIT=16'h0100;
LUT4 \top/uart_rx_inst/state_0_s6  (
	.I0(\top/uart_rx_inst/bit_cnt [3]),
	.I1(\top/uart_rx_inst/bit_cnt [1]),
	.I2(\top/uart_rx_inst/bit_cnt [2]),
	.I3(\top/uart_rx_inst/bit_cnt [0]),
	.F(\top/uart_rx_inst/state_0_11 )
);
defparam \top/uart_rx_inst/state_0_s6 .INIT=16'h4000;
LUT4 \top/uart_rx_inst/rx_data_7_s3  (
	.I0(rst),
	.I1(\top/uart_rx_inst/state [0]),
	.I2(\top/uart_rx_inst/state [1]),
	.I3(\top/uart_rx_inst/n191_10 ),
	.F(\top/uart_rx_inst/rx_data_7_6 )
);
defparam \top/uart_rx_inst/rx_data_7_s3 .INIT=16'h4000;
LUT4 \top/uart_rx_inst/shift_reg_7_s5  (
	.I0(rst),
	.I1(\top/uart_rx_inst/state [0]),
	.I2(\top/uart_rx_inst/state [1]),
	.I3(\top/uart_rx_inst/n191_10 ),
	.F(\top/uart_rx_inst/shift_reg_7_10 )
);
defparam \top/uart_rx_inst/shift_reg_7_s5 .INIT=16'h1400;
LUT4 \top/uart_rx_inst/n217_s8  (
	.I0(\top/uart_rx_inst/n191_10 ),
	.I1(\top/uart_rx_inst/rx_dd ),
	.I2(\top/uart_rx_inst/state [0]),
	.I3(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/n217_14 )
);
defparam \top/uart_rx_inst/n217_s8 .INIT=16'h555C;
LUT4 \top/uart_rx_inst/n22_s3  (
	.I0(\top/uart_rx_inst/state [0]),
	.I1(\top/uart_rx_inst/state [1]),
	.I2(\top/uart_rx_inst/baud_cnt [1]),
	.I3(\top/uart_rx_inst/baud_cnt [0]),
	.F(\top/uart_rx_inst/n22_8 )
);
defparam \top/uart_rx_inst/n22_s3 .INIT=16'h1FF1;
LUT3 \top/uart_rx_inst/baud_cnt_8_s3  (
	.I0(\top/uart_rx_inst/rx_dd ),
	.I1(\top/uart_rx_inst/state [0]),
	.I2(\top/uart_rx_inst/state [1]),
	.F(\top/uart_rx_inst/baud_cnt_8_9 )
);
defparam \top/uart_rx_inst/baud_cnt_8_s3 .INIT=8'hFD;
DFFC \top/uart_rx_inst/rx_valid_s0  (
	.D(\top/uart_rx_inst/n191_9 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/rx_valid_Z )
);
defparam \top/uart_rx_inst/rx_valid_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_d_s0  (
	.D(uart_rx),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_d_7 ),
	.Q(\top/uart_rx_inst/rx_d )
);
defparam \top/uart_rx_inst/rx_d_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_dd_s0  (
	.D(\top/uart_rx_inst/rx_d ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_d_7 ),
	.Q(\top/uart_rx_inst/rx_dd )
);
defparam \top/uart_rx_inst/rx_dd_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_7_s0  (
	.D(\top/uart_rx_inst/shift_reg [7]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [7])
);
defparam \top/uart_rx_inst/rx_data_7_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_6_s0  (
	.D(\top/uart_rx_inst/shift_reg [6]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [6])
);
defparam \top/uart_rx_inst/rx_data_6_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_5_s0  (
	.D(\top/uart_rx_inst/shift_reg [5]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [5])
);
defparam \top/uart_rx_inst/rx_data_5_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_4_s0  (
	.D(\top/uart_rx_inst/shift_reg [4]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [4])
);
defparam \top/uart_rx_inst/rx_data_4_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_3_s0  (
	.D(\top/uart_rx_inst/shift_reg [3]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [3])
);
defparam \top/uart_rx_inst/rx_data_3_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_2_s0  (
	.D(\top/uart_rx_inst/shift_reg [2]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [2])
);
defparam \top/uart_rx_inst/rx_data_2_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_1_s0  (
	.D(\top/uart_rx_inst/shift_reg [1]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [1])
);
defparam \top/uart_rx_inst/rx_data_1_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/rx_data_0_s0  (
	.D(\top/uart_rx_inst/shift_reg [0]),
	.CLK(clk),
	.CE(\top/uart_rx_inst/rx_data_7_6 ),
	.Q(\top/rx_data_Z [0])
);
defparam \top/uart_rx_inst/rx_data_0_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_7_s0  (
	.D(\top/uart_rx_inst/n218_12 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [7])
);
defparam \top/uart_rx_inst/shift_reg_7_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_6_s0  (
	.D(\top/uart_rx_inst/n219_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [6])
);
defparam \top/uart_rx_inst/shift_reg_6_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_5_s0  (
	.D(\top/uart_rx_inst/n220_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [5])
);
defparam \top/uart_rx_inst/shift_reg_5_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_4_s0  (
	.D(\top/uart_rx_inst/n221_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [4])
);
defparam \top/uart_rx_inst/shift_reg_4_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_3_s0  (
	.D(\top/uart_rx_inst/n222_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [3])
);
defparam \top/uart_rx_inst/shift_reg_3_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_2_s0  (
	.D(\top/uart_rx_inst/n223_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [2])
);
defparam \top/uart_rx_inst/shift_reg_2_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_1_s0  (
	.D(\top/uart_rx_inst/n224_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [1])
);
defparam \top/uart_rx_inst/shift_reg_1_s0 .INIT=1'b0;
DFFE \top/uart_rx_inst/shift_reg_0_s0  (
	.D(\top/uart_rx_inst/n225_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/shift_reg_7_10 ),
	.Q(\top/uart_rx_inst/shift_reg [0])
);
defparam \top/uart_rx_inst/shift_reg_0_s0 .INIT=1'b0;
DFFCE \top/uart_rx_inst/bit_cnt_3_s1  (
	.D(\top/uart_rx_inst/n226_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/bit_cnt_3_8 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/bit_cnt [3])
);
defparam \top/uart_rx_inst/bit_cnt_3_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/bit_cnt_2_s1  (
	.D(\top/uart_rx_inst/n227_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/bit_cnt_3_8 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/bit_cnt [2])
);
defparam \top/uart_rx_inst/bit_cnt_2_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/bit_cnt_1_s1  (
	.D(\top/uart_rx_inst/n228_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/bit_cnt_3_8 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/bit_cnt [1])
);
defparam \top/uart_rx_inst/bit_cnt_1_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/bit_cnt_0_s1  (
	.D(\top/uart_rx_inst/n229_12 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/bit_cnt_3_8 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/bit_cnt [0])
);
defparam \top/uart_rx_inst/bit_cnt_0_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_15_s1  (
	.D(\top/uart_rx_inst/n202_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [15])
);
defparam \top/uart_rx_inst/baud_cnt_15_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_14_s1  (
	.D(\top/uart_rx_inst/n203_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [14])
);
defparam \top/uart_rx_inst/baud_cnt_14_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_13_s1  (
	.D(\top/uart_rx_inst/n204_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [13])
);
defparam \top/uart_rx_inst/baud_cnt_13_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_12_s1  (
	.D(\top/uart_rx_inst/n205_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [12])
);
defparam \top/uart_rx_inst/baud_cnt_12_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_11_s1  (
	.D(\top/uart_rx_inst/n206_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [11])
);
defparam \top/uart_rx_inst/baud_cnt_11_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_10_s1  (
	.D(\top/uart_rx_inst/n207_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [10])
);
defparam \top/uart_rx_inst/baud_cnt_10_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_9_s1  (
	.D(\top/uart_rx_inst/n208_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [9])
);
defparam \top/uart_rx_inst/baud_cnt_9_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_8_s1  (
	.D(\top/uart_rx_inst/n15_6 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [8])
);
defparam \top/uart_rx_inst/baud_cnt_8_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_7_s1  (
	.D(\top/uart_rx_inst/n16_6 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [7])
);
defparam \top/uart_rx_inst/baud_cnt_7_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_6_s1  (
	.D(\top/uart_rx_inst/n211_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [6])
);
defparam \top/uart_rx_inst/baud_cnt_6_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_5_s1  (
	.D(\top/uart_rx_inst/n18_6 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [5])
);
defparam \top/uart_rx_inst/baud_cnt_5_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_4_s1  (
	.D(\top/uart_rx_inst/n19_6 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [4])
);
defparam \top/uart_rx_inst/baud_cnt_4_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_3_s1  (
	.D(\top/uart_rx_inst/n214_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [3])
);
defparam \top/uart_rx_inst/baud_cnt_3_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_2_s1  (
	.D(\top/uart_rx_inst/n215_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [2])
);
defparam \top/uart_rx_inst/baud_cnt_2_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_1_s1  (
	.D(\top/uart_rx_inst/n22_8 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [1])
);
defparam \top/uart_rx_inst/baud_cnt_1_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/baud_cnt_0_s1  (
	.D(\top/uart_rx_inst/n217_11 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/baud_cnt_8_9 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/baud_cnt [0])
);
defparam \top/uart_rx_inst/baud_cnt_0_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/state_1_s1  (
	.D(\top/uart_rx_inst/n200_12 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/n139_4 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/state [1])
);
defparam \top/uart_rx_inst/state_1_s1 .INIT=1'b0;
DFFCE \top/uart_rx_inst/state_0_s1  (
	.D(\top/uart_rx_inst/n201_20 ),
	.CLK(clk),
	.CE(\top/uart_rx_inst/n139_4 ),
	.CLEAR(rst),
	.Q(\top/uart_rx_inst/state [0])
);
defparam \top/uart_rx_inst/state_0_s1 .INIT=1'b0;
INV \top/uart_rx_inst/rx_d_s3  (
	.I(rst),
	.O(\top/uart_rx_inst/rx_d_7 )
);
LUT1 \top/uart_rx_inst/n201_s14  (
	.I0(\top/uart_rx_inst/state [0]),
	.F(\top/uart_rx_inst/n201_20 )
);
defparam \top/uart_rx_inst/n201_s14 .INIT=2'h1;
LUT4 \top/uart_tx_inst/tx_s3  (
	.I0(\top/uart_tx_inst/tx_6 ),
	.I1(\top/uart_tx_inst/baud_cnt [8]),
	.I2(\top/uart_tx_inst/baud_cnt [9]),
	.I3(\top/uart_tx_inst/tx_7 ),
	.F(\top/uart_tx_inst/tx_5 )
);
defparam \top/uart_tx_inst/tx_s3 .INIT=16'h40FF;
LUT2 \top/uart_tx_inst/n113_s6  (
	.I0(\top/uart_tx_inst/baud_cnt [0]),
	.I1(\top/uart_tx_inst/n80_7 ),
	.F(\top/uart_tx_inst/n113_11 )
);
defparam \top/uart_tx_inst/n113_s6 .INIT=4'h1;
LUT3 \top/uart_tx_inst/n112_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [1]),
	.I2(\top/uart_tx_inst/baud_cnt [0]),
	.F(\top/uart_tx_inst/n112_11 )
);
defparam \top/uart_tx_inst/n112_s6 .INIT=8'h14;
LUT4 \top/uart_tx_inst/n110_s6  (
	.I0(\top/uart_tx_inst/baud_cnt [2]),
	.I1(\top/uart_tx_inst/n111_12 ),
	.I2(\top/uart_tx_inst/n80_7 ),
	.I3(\top/uart_tx_inst/baud_cnt [3]),
	.F(\top/uart_tx_inst/n110_11 )
);
defparam \top/uart_tx_inst/n110_s6 .INIT=16'h0708;
LUT3 \top/uart_tx_inst/n109_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [4]),
	.I2(\top/uart_tx_inst/n109_14 ),
	.F(\top/uart_tx_inst/n109_11 )
);
defparam \top/uart_tx_inst/n109_s6 .INIT=8'h14;
LUT4 \top/uart_tx_inst/n108_s6  (
	.I0(\top/uart_tx_inst/baud_cnt [4]),
	.I1(\top/uart_tx_inst/n109_14 ),
	.I2(\top/uart_tx_inst/n80_7 ),
	.I3(\top/uart_tx_inst/baud_cnt [5]),
	.F(\top/uart_tx_inst/n108_11 )
);
defparam \top/uart_tx_inst/n108_s6 .INIT=16'h0708;
LUT3 \top/uart_tx_inst/n107_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/n107_12 ),
	.I2(\top/uart_tx_inst/baud_cnt [6]),
	.F(\top/uart_tx_inst/n107_11 )
);
defparam \top/uart_tx_inst/n107_s6 .INIT=8'h14;
LUT3 \top/uart_tx_inst/n106_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [7]),
	.I2(\top/uart_tx_inst/n106_12 ),
	.F(\top/uart_tx_inst/n106_11 )
);
defparam \top/uart_tx_inst/n106_s6 .INIT=8'h14;
LUT4 \top/uart_tx_inst/n104_s6  (
	.I0(\top/uart_tx_inst/baud_cnt [8]),
	.I1(\top/uart_tx_inst/n105_12 ),
	.I2(\top/uart_tx_inst/n80_7 ),
	.I3(\top/uart_tx_inst/baud_cnt [9]),
	.F(\top/uart_tx_inst/n104_11 )
);
defparam \top/uart_tx_inst/n104_s6 .INIT=16'h0708;
LUT3 \top/uart_tx_inst/n103_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/n103_14 ),
	.I2(\top/uart_tx_inst/baud_cnt [10]),
	.F(\top/uart_tx_inst/n103_11 )
);
defparam \top/uart_tx_inst/n103_s6 .INIT=8'h14;
LUT3 \top/uart_tx_inst/n102_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [11]),
	.I2(\top/uart_tx_inst/n102_12 ),
	.F(\top/uart_tx_inst/n102_11 )
);
defparam \top/uart_tx_inst/n102_s6 .INIT=8'h14;
LUT4 \top/uart_tx_inst/n101_s6  (
	.I0(\top/uart_tx_inst/baud_cnt [11]),
	.I1(\top/uart_tx_inst/n102_12 ),
	.I2(\top/uart_tx_inst/n80_7 ),
	.I3(\top/uart_tx_inst/baud_cnt [12]),
	.F(\top/uart_tx_inst/n101_11 )
);
defparam \top/uart_tx_inst/n101_s6 .INIT=16'h0708;
LUT3 \top/uart_tx_inst/n100_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/n100_12 ),
	.I2(\top/uart_tx_inst/baud_cnt [13]),
	.F(\top/uart_tx_inst/n100_11 )
);
defparam \top/uart_tx_inst/n100_s6 .INIT=8'h14;
LUT3 \top/uart_tx_inst/n99_s6  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [14]),
	.I2(\top/uart_tx_inst/n99_12 ),
	.F(\top/uart_tx_inst/n99_11 )
);
defparam \top/uart_tx_inst/n99_s6 .INIT=8'h14;
LUT4 \top/uart_tx_inst/n98_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [14]),
	.I1(\top/uart_tx_inst/n99_12 ),
	.I2(\top/uart_tx_inst/n80_7 ),
	.I3(\top/uart_tx_inst/baud_cnt [15]),
	.F(\top/uart_tx_inst/n98_13 )
);
defparam \top/uart_tx_inst/n98_s7 .INIT=16'h0708;
LUT4 \top/uart_tx_inst/n126_s5  (
	.I0(\top/uart_tx_inst/bit_index [0]),
	.I1(\top/uart_tx_inst/bit_index [1]),
	.I2(\top/uart_tx_inst/tx_busy_9 ),
	.I3(\top/uart_tx_inst/bit_index [2]),
	.F(\top/uart_tx_inst/n126_10 )
);
defparam \top/uart_tx_inst/n126_s5 .INIT=16'h0708;
LUT4 \top/uart_tx_inst/tx_s4  (
	.I0(\top/uart_tx_inst/tx_8 ),
	.I1(\top/uart_tx_inst/baud_cnt [6]),
	.I2(\top/uart_tx_inst/baud_cnt [5]),
	.I3(\top/uart_tx_inst/baud_cnt [7]),
	.F(\top/uart_tx_inst/tx_6 )
);
defparam \top/uart_tx_inst/tx_s4 .INIT=16'h00BF;
LUT4 \top/uart_tx_inst/tx_s5  (
	.I0(\top/uart_tx_inst/baud_cnt [10]),
	.I1(\top/uart_tx_inst/baud_cnt [11]),
	.I2(\top/uart_tx_inst/tx_busy_9 ),
	.I3(\top/uart_tx_inst/tx_9 ),
	.F(\top/uart_tx_inst/tx_7 )
);
defparam \top/uart_tx_inst/tx_s5 .INIT=16'h0100;
LUT2 \top/uart_tx_inst/n111_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [1]),
	.I1(\top/uart_tx_inst/baud_cnt [0]),
	.F(\top/uart_tx_inst/n111_12 )
);
defparam \top/uart_tx_inst/n111_s7 .INIT=4'h8;
LUT3 \top/uart_tx_inst/n107_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [4]),
	.I1(\top/uart_tx_inst/baud_cnt [5]),
	.I2(\top/uart_tx_inst/n109_14 ),
	.F(\top/uart_tx_inst/n107_12 )
);
defparam \top/uart_tx_inst/n107_s7 .INIT=8'h80;
LUT4 \top/uart_tx_inst/n106_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [4]),
	.I1(\top/uart_tx_inst/baud_cnt [5]),
	.I2(\top/uart_tx_inst/baud_cnt [6]),
	.I3(\top/uart_tx_inst/n109_14 ),
	.F(\top/uart_tx_inst/n106_12 )
);
defparam \top/uart_tx_inst/n106_s7 .INIT=16'h8000;
LUT2 \top/uart_tx_inst/n105_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [7]),
	.I1(\top/uart_tx_inst/n106_12 ),
	.F(\top/uart_tx_inst/n105_12 )
);
defparam \top/uart_tx_inst/n105_s7 .INIT=4'h8;
LUT4 \top/uart_tx_inst/n102_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [8]),
	.I1(\top/uart_tx_inst/baud_cnt [9]),
	.I2(\top/uart_tx_inst/baud_cnt [10]),
	.I3(\top/uart_tx_inst/n105_12 ),
	.F(\top/uart_tx_inst/n102_12 )
);
defparam \top/uart_tx_inst/n102_s7 .INIT=16'h8000;
LUT3 \top/uart_tx_inst/n100_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [11]),
	.I1(\top/uart_tx_inst/baud_cnt [12]),
	.I2(\top/uart_tx_inst/n102_12 ),
	.F(\top/uart_tx_inst/n100_12 )
);
defparam \top/uart_tx_inst/n100_s7 .INIT=8'h80;
LUT4 \top/uart_tx_inst/n99_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [11]),
	.I1(\top/uart_tx_inst/baud_cnt [12]),
	.I2(\top/uart_tx_inst/baud_cnt [13]),
	.I3(\top/uart_tx_inst/n102_12 ),
	.F(\top/uart_tx_inst/n99_12 )
);
defparam \top/uart_tx_inst/n99_s7 .INIT=16'h8000;
LUT4 \top/uart_tx_inst/n129_s6  (
	.I0(\top/uart_tx_inst/bit_index [1]),
	.I1(\top/uart_tx_inst/bit_index [2]),
	.I2(\top/uart_tx_inst/bit_index [0]),
	.I3(\top/uart_tx_inst/bit_index [3]),
	.F(\top/uart_tx_inst/n129_11 )
);
defparam \top/uart_tx_inst/n129_s6 .INIT=16'h1000;
LUT3 \top/uart_tx_inst/n125_s6  (
	.I0(\top/uart_tx_inst/bit_index [0]),
	.I1(\top/uart_tx_inst/bit_index [1]),
	.I2(\top/uart_tx_inst/bit_index [2]),
	.F(\top/uart_tx_inst/n125_11 )
);
defparam \top/uart_tx_inst/n125_s6 .INIT=8'h80;
LUT4 \top/uart_tx_inst/tx_s6  (
	.I0(\top/uart_tx_inst/baud_cnt [2]),
	.I1(\top/uart_tx_inst/baud_cnt [3]),
	.I2(\top/uart_tx_inst/baud_cnt [4]),
	.I3(\top/uart_tx_inst/n111_12 ),
	.F(\top/uart_tx_inst/tx_8 )
);
defparam \top/uart_tx_inst/tx_s6 .INIT=16'h0001;
LUT4 \top/uart_tx_inst/tx_s7  (
	.I0(\top/uart_tx_inst/baud_cnt [12]),
	.I1(\top/uart_tx_inst/baud_cnt [13]),
	.I2(\top/uart_tx_inst/baud_cnt [14]),
	.I3(\top/uart_tx_inst/baud_cnt [15]),
	.F(\top/uart_tx_inst/tx_9 )
);
defparam \top/uart_tx_inst/tx_s7 .INIT=16'h0001;
LUT4 \top/uart_tx_inst/n103_s8  (
	.I0(\top/uart_tx_inst/baud_cnt [8]),
	.I1(\top/uart_tx_inst/baud_cnt [9]),
	.I2(\top/uart_tx_inst/baud_cnt [7]),
	.I3(\top/uart_tx_inst/n106_12 ),
	.F(\top/uart_tx_inst/n103_14 )
);
defparam \top/uart_tx_inst/n103_s8 .INIT=16'h8000;
LUT4 \top/uart_tx_inst/n105_s8  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [8]),
	.I2(\top/uart_tx_inst/baud_cnt [7]),
	.I3(\top/uart_tx_inst/n106_12 ),
	.F(\top/uart_tx_inst/n105_14 )
);
defparam \top/uart_tx_inst/n105_s8 .INIT=16'h1444;
LUT4 \top/uart_tx_inst/n109_s8  (
	.I0(\top/uart_tx_inst/baud_cnt [2]),
	.I1(\top/uart_tx_inst/baud_cnt [3]),
	.I2(\top/uart_tx_inst/baud_cnt [1]),
	.I3(\top/uart_tx_inst/baud_cnt [0]),
	.F(\top/uart_tx_inst/n109_14 )
);
defparam \top/uart_tx_inst/n109_s8 .INIT=16'h8000;
LUT4 \top/uart_tx_inst/n111_s8  (
	.I0(\top/uart_tx_inst/n80_7 ),
	.I1(\top/uart_tx_inst/baud_cnt [2]),
	.I2(\top/uart_tx_inst/baud_cnt [1]),
	.I3(\top/uart_tx_inst/baud_cnt [0]),
	.F(\top/uart_tx_inst/n111_14 )
);
defparam \top/uart_tx_inst/n111_s8 .INIT=16'h1444;
LUT3 \top/uart_tx_inst/n81_s3  (
	.I0(\top/uart_tx_inst/shift_reg [0]),
	.I1(\top/uart_tx_inst/state [0]),
	.I2(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n81_8 )
);
defparam \top/uart_tx_inst/n81_s3 .INIT=8'hAB;
LUT3 \top/uart_tx_inst/n124_s6  (
	.I0(\top/uart_tx_inst/state [0]),
	.I1(\top/uart_tx_inst/state [1]),
	.I2(\top/uart_tx_inst/shift_reg [1]),
	.F(\top/uart_tx_inst/n124_12 )
);
defparam \top/uart_tx_inst/n124_s6 .INIT=8'hE0;
LUT4 \top/uart_tx_inst/n125_s7  (
	.I0(\top/uart_tx_inst/state [0]),
	.I1(\top/uart_tx_inst/state [1]),
	.I2(\top/uart_tx_inst/n125_11 ),
	.I3(\top/uart_tx_inst/bit_index [3]),
	.F(\top/uart_tx_inst/n125_13 )
);
defparam \top/uart_tx_inst/n125_s7 .INIT=16'h0EE0;
LUT4 \top/uart_tx_inst/n127_s6  (
	.I0(\top/uart_tx_inst/state [0]),
	.I1(\top/uart_tx_inst/state [1]),
	.I2(\top/uart_tx_inst/bit_index [0]),
	.I3(\top/uart_tx_inst/bit_index [1]),
	.F(\top/uart_tx_inst/n127_12 )
);
defparam \top/uart_tx_inst/n127_s6 .INIT=16'h0EE0;
LUT3 \top/uart_tx_inst/n128_s7  (
	.I0(\top/uart_tx_inst/bit_index [0]),
	.I1(\top/uart_tx_inst/state [0]),
	.I2(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n128_13 )
);
defparam \top/uart_tx_inst/n128_s7 .INIT=8'h54;
LUT3 \top/uart_tx_inst/n129_s7  (
	.I0(\top/uart_tx_inst/n129_11 ),
	.I1(\top/uart_tx_inst/state [0]),
	.I2(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n129_13 )
);
defparam \top/uart_tx_inst/n129_s7 .INIT=8'h54;
LUT3 \top/uart_tx_inst/baud_cnt_15_s4  (
	.I0(\top/tx_start ),
	.I1(\top/uart_tx_inst/state [0]),
	.I2(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/baud_cnt_15_10 )
);
defparam \top/uart_tx_inst/baud_cnt_15_s4 .INIT=8'hFE;
LUT2 \top/uart_tx_inst/n98_s8  (
	.I0(\top/uart_tx_inst/state [0]),
	.I1(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n98_15 )
);
defparam \top/uart_tx_inst/n98_s8 .INIT=4'hE;
LUT4 \top/uart_tx_inst/n123_s5  (
	.I0(\top/uart_tx_inst/shift_reg [2]),
	.I1(\top/tx_data [0]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n123_10 )
);
defparam \top/uart_tx_inst/n123_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/n122_s5  (
	.I0(\top/uart_tx_inst/shift_reg [3]),
	.I1(\top/tx_data [1]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n122_10 )
);
defparam \top/uart_tx_inst/n122_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/n121_s5  (
	.I0(\top/uart_tx_inst/shift_reg [4]),
	.I1(\top/tx_data [2]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n121_10 )
);
defparam \top/uart_tx_inst/n121_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/n120_s5  (
	.I0(\top/uart_tx_inst/shift_reg [5]),
	.I1(\top/tx_data [3]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n120_10 )
);
defparam \top/uart_tx_inst/n120_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/n119_s5  (
	.I0(\top/uart_tx_inst/shift_reg [6]),
	.I1(\top/tx_data [4]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n119_10 )
);
defparam \top/uart_tx_inst/n119_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/n118_s5  (
	.I0(\top/uart_tx_inst/shift_reg [7]),
	.I1(\top/tx_data [5]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n118_10 )
);
defparam \top/uart_tx_inst/n118_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/n117_s5  (
	.I0(\top/uart_tx_inst/shift_reg [8]),
	.I1(\top/tx_data [6]),
	.I2(\top/uart_tx_inst/state [0]),
	.I3(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/n117_10 )
);
defparam \top/uart_tx_inst/n117_s5 .INIT=16'hAAAC;
LUT4 \top/uart_tx_inst/tx_busy_s4  (
	.I0(\top/uart_tx_inst/state [0]),
	.I1(\top/uart_tx_inst/state [1]),
	.I2(\top/uart_tx_inst/baud_cnt_15_10 ),
	.I3(\top/uart_tx_inst/tx_5 ),
	.F(\top/uart_tx_inst/tx_busy_7 )
);
defparam \top/uart_tx_inst/tx_busy_s4 .INIT=16'h1AAA;
LUT2 \top/uart_tx_inst/tx_busy_s5  (
	.I0(\top/uart_tx_inst/state [0]),
	.I1(\top/uart_tx_inst/state [1]),
	.F(\top/uart_tx_inst/tx_busy_9 )
);
defparam \top/uart_tx_inst/tx_busy_s5 .INIT=4'h1;
LUT4 \top/uart_tx_inst/n80_s2  (
	.I0(\top/tx_start ),
	.I1(\top/uart_tx_inst/state [0]),
	.I2(\top/uart_tx_inst/state [1]),
	.I3(\top/uart_tx_inst/tx_5 ),
	.F(\top/uart_tx_inst/n80_7 )
);
defparam \top/uart_tx_inst/n80_s2 .INIT=16'hFE00;
DFFCE \top/uart_tx_inst/tx_busy_s0  (
	.D(\top/tx_start ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/tx_busy_9 ),
	.CLEAR(rst),
	.Q(\top/tx_busy_Z )
);
defparam \top/uart_tx_inst/tx_busy_s0 .INIT=1'b0;
DFFCE \top/uart_tx_inst/state_1_s1  (
	.D(\top/uart_tx_inst/n129_13 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/state [1])
);
defparam \top/uart_tx_inst/state_1_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_15_s1  (
	.D(\top/uart_tx_inst/n98_13 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [15])
);
defparam \top/uart_tx_inst/baud_cnt_15_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_14_s1  (
	.D(\top/uart_tx_inst/n99_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [14])
);
defparam \top/uart_tx_inst/baud_cnt_14_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_13_s1  (
	.D(\top/uart_tx_inst/n100_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [13])
);
defparam \top/uart_tx_inst/baud_cnt_13_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_12_s1  (
	.D(\top/uart_tx_inst/n101_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [12])
);
defparam \top/uart_tx_inst/baud_cnt_12_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_11_s1  (
	.D(\top/uart_tx_inst/n102_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [11])
);
defparam \top/uart_tx_inst/baud_cnt_11_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_10_s1  (
	.D(\top/uart_tx_inst/n103_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [10])
);
defparam \top/uart_tx_inst/baud_cnt_10_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_9_s1  (
	.D(\top/uart_tx_inst/n104_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [9])
);
defparam \top/uart_tx_inst/baud_cnt_9_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_8_s1  (
	.D(\top/uart_tx_inst/n105_14 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [8])
);
defparam \top/uart_tx_inst/baud_cnt_8_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_7_s1  (
	.D(\top/uart_tx_inst/n106_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [7])
);
defparam \top/uart_tx_inst/baud_cnt_7_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_6_s1  (
	.D(\top/uart_tx_inst/n107_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [6])
);
defparam \top/uart_tx_inst/baud_cnt_6_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_5_s1  (
	.D(\top/uart_tx_inst/n108_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [5])
);
defparam \top/uart_tx_inst/baud_cnt_5_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_4_s1  (
	.D(\top/uart_tx_inst/n109_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [4])
);
defparam \top/uart_tx_inst/baud_cnt_4_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_3_s1  (
	.D(\top/uart_tx_inst/n110_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [3])
);
defparam \top/uart_tx_inst/baud_cnt_3_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_2_s1  (
	.D(\top/uart_tx_inst/n111_14 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [2])
);
defparam \top/uart_tx_inst/baud_cnt_2_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_1_s1  (
	.D(\top/uart_tx_inst/n112_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [1])
);
defparam \top/uart_tx_inst/baud_cnt_1_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/baud_cnt_0_s1  (
	.D(\top/uart_tx_inst/n113_11 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/baud_cnt_15_10 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/baud_cnt [0])
);
defparam \top/uart_tx_inst/baud_cnt_0_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/bit_index_3_s1  (
	.D(\top/uart_tx_inst/n125_13 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/bit_index [3])
);
defparam \top/uart_tx_inst/bit_index_3_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/bit_index_2_s1  (
	.D(\top/uart_tx_inst/n126_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/bit_index [2])
);
defparam \top/uart_tx_inst/bit_index_2_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/bit_index_1_s1  (
	.D(\top/uart_tx_inst/n127_12 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/bit_index [1])
);
defparam \top/uart_tx_inst/bit_index_1_s1 .INIT=1'b0;
DFFCE \top/uart_tx_inst/bit_index_0_s1  (
	.D(\top/uart_tx_inst/n128_13 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/bit_index [0])
);
defparam \top/uart_tx_inst/bit_index_0_s1 .INIT=1'b0;
DFFPE \top/uart_tx_inst/shift_reg_8_s1  (
	.D(\top/uart_tx_inst/n98_15 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [8])
);
defparam \top/uart_tx_inst/shift_reg_8_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_7_s1  (
	.D(\top/uart_tx_inst/n117_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [7])
);
defparam \top/uart_tx_inst/shift_reg_7_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_6_s1  (
	.D(\top/uart_tx_inst/n118_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [6])
);
defparam \top/uart_tx_inst/shift_reg_6_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_5_s1  (
	.D(\top/uart_tx_inst/n119_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [5])
);
defparam \top/uart_tx_inst/shift_reg_5_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_4_s1  (
	.D(\top/uart_tx_inst/n120_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [4])
);
defparam \top/uart_tx_inst/shift_reg_4_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_3_s1  (
	.D(\top/uart_tx_inst/n121_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [3])
);
defparam \top/uart_tx_inst/shift_reg_3_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_2_s1  (
	.D(\top/uart_tx_inst/n122_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [2])
);
defparam \top/uart_tx_inst/shift_reg_2_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_1_s1  (
	.D(\top/uart_tx_inst/n123_10 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [1])
);
defparam \top/uart_tx_inst/shift_reg_1_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/shift_reg_0_s1  (
	.D(\top/uart_tx_inst/n124_12 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/n80_7 ),
	.PRESET(rst),
	.Q(\top/uart_tx_inst/shift_reg [0])
);
defparam \top/uart_tx_inst/shift_reg_0_s1 .INIT=1'b1;
DFFPE \top/uart_tx_inst/tx_s1  (
	.D(\top/uart_tx_inst/n81_8 ),
	.CLK(clk),
	.CE(\top/uart_tx_inst/tx_5 ),
	.PRESET(rst),
	.Q(uart_tx)
);
defparam \top/uart_tx_inst/tx_s1 .INIT=1'b1;
DFFC \top/uart_tx_inst/state_0_s2  (
	.D(\top/uart_tx_inst/tx_busy_7 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/uart_tx_inst/state [0])
);
defparam \top/uart_tx_inst/state_0_s2 .INIT=1'b0;
LUT3 \top/processor/n7631_s0  (
	.I0(\top/processor/n7631_8 ),
	.I1(\top/processor/n7631_12 ),
	.I2(\top/processor/n7631_10 ),
	.F(\top/processor/n7631_3 )
);
defparam \top/processor/n7631_s0 .INIT=8'h8F;
LUT4 \top/processor/n10817_s9  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/n10817_15 ),
	.I2(\top/data_in [7]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n10817_14 )
);
defparam \top/processor/n10817_s9 .INIT=16'hEEF0;
LUT4 \top/processor/n10825_s9  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/n10817_15 ),
	.I2(\top/data_in [7]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n10825_14 )
);
defparam \top/processor/n10825_s9 .INIT=16'h44F0;
LUT4 \top/processor/n11265_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [63]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11265_12 )
);
defparam \top/processor/n11265_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11266_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [62]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11266_12 )
);
defparam \top/processor/n11266_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11267_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [61]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11267_12 )
);
defparam \top/processor/n11267_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11268_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [60]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11268_12 )
);
defparam \top/processor/n11268_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11269_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [59]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11269_12 )
);
defparam \top/processor/n11269_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11270_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [58]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11270_12 )
);
defparam \top/processor/n11270_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11271_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [57]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11271_12 )
);
defparam \top/processor/n11271_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11272_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [56]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11272_12 )
);
defparam \top/processor/n11272_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11273_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [55]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11273_12 )
);
defparam \top/processor/n11273_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11274_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [54]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11274_12 )
);
defparam \top/processor/n11274_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11275_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [53]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11275_12 )
);
defparam \top/processor/n11275_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11276_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [52]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11276_12 )
);
defparam \top/processor/n11276_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11277_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [51]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11277_12 )
);
defparam \top/processor/n11277_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11278_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [50]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11278_12 )
);
defparam \top/processor/n11278_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11279_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [49]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11279_12 )
);
defparam \top/processor/n11279_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11280_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [48]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11280_12 )
);
defparam \top/processor/n11280_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11281_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [47]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11281_12 )
);
defparam \top/processor/n11281_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11282_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [46]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11282_12 )
);
defparam \top/processor/n11282_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11283_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [45]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11283_12 )
);
defparam \top/processor/n11283_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11284_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [44]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11284_12 )
);
defparam \top/processor/n11284_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11285_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [43]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11285_12 )
);
defparam \top/processor/n11285_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11286_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [42]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11286_12 )
);
defparam \top/processor/n11286_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11287_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [41]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11287_12 )
);
defparam \top/processor/n11287_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11288_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [40]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11288_12 )
);
defparam \top/processor/n11288_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11289_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [39]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11289_12 )
);
defparam \top/processor/n11289_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11290_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [38]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11290_12 )
);
defparam \top/processor/n11290_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11291_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [37]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11291_12 )
);
defparam \top/processor/n11291_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11292_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [36]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11292_12 )
);
defparam \top/processor/n11292_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11293_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [35]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11293_12 )
);
defparam \top/processor/n11293_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11294_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [34]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11294_12 )
);
defparam \top/processor/n11294_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11295_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [33]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11295_12 )
);
defparam \top/processor/n11295_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11296_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [32]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11296_12 )
);
defparam \top/processor/n11296_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11297_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [31]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11297_12 )
);
defparam \top/processor/n11297_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11298_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [30]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11298_12 )
);
defparam \top/processor/n11298_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11299_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [29]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11299_12 )
);
defparam \top/processor/n11299_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11300_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [28]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11300_12 )
);
defparam \top/processor/n11300_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11301_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [27]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11301_12 )
);
defparam \top/processor/n11301_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11302_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [26]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11302_12 )
);
defparam \top/processor/n11302_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11303_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [25]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11303_12 )
);
defparam \top/processor/n11303_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11304_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [24]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11304_12 )
);
defparam \top/processor/n11304_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11305_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [23]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11305_12 )
);
defparam \top/processor/n11305_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11306_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [22]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11306_12 )
);
defparam \top/processor/n11306_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11307_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [21]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11307_12 )
);
defparam \top/processor/n11307_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11308_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [20]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11308_12 )
);
defparam \top/processor/n11308_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11309_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [19]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11309_12 )
);
defparam \top/processor/n11309_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11310_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [18]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11310_12 )
);
defparam \top/processor/n11310_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11311_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [17]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11311_12 )
);
defparam \top/processor/n11311_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11312_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [16]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11312_12 )
);
defparam \top/processor/n11312_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11313_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [15]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11313_12 )
);
defparam \top/processor/n11313_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11314_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [14]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11314_12 )
);
defparam \top/processor/n11314_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11315_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [13]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11315_12 )
);
defparam \top/processor/n11315_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11316_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [12]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11316_12 )
);
defparam \top/processor/n11316_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11317_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [11]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11317_12 )
);
defparam \top/processor/n11317_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11318_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [10]),
	.I2(\top/data_in [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11318_12 )
);
defparam \top/processor/n11318_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11319_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [9]),
	.I2(\top/data_in [1]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11319_12 )
);
defparam \top/processor/n11319_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11320_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [8]),
	.I2(\top/data_in [0]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11320_12 )
);
defparam \top/processor/n11320_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11321_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/total_bits [7]),
	.I3(\top/processor/n10825_14 ),
	.F(\top/processor/n11321_12 )
);
defparam \top/processor/n11321_s8 .INIT=16'hFF40;
LUT4 \top/processor/n11322_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [6]),
	.I2(\top/data_in [6]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11322_12 )
);
defparam \top/processor/n11322_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11323_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [5]),
	.I2(\top/data_in [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11323_12 )
);
defparam \top/processor/n11323_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11324_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [4]),
	.I2(\top/data_in [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11324_12 )
);
defparam \top/processor/n11324_s8 .INIT=16'h44F0;
LUT4 \top/processor/n11325_s8  (
	.I0(\top/processor/n11265_13 ),
	.I1(\top/processor/total_bits [3]),
	.I2(\top/data_in [3]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11325_12 )
);
defparam \top/processor/n11325_s8 .INIT=16'h44F0;
LUT3 \top/processor/n11361_s10  (
	.I0(\top/processor/n11361_17 ),
	.I1(\top/state_0 [0]),
	.I2(\top/state_0 [1]),
	.F(\top/processor/n11361_16 )
);
defparam \top/processor/n11361_s10 .INIT=8'h2C;
LUT2 \top/processor/n11363_s10  (
	.I0(\top/state_0 [0]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n11363_16 )
);
defparam \top/processor/n11363_s10 .INIT=4'h6;
LUT4 \top/processor/n11364_s21  (
	.I0(\top/processor/need_length_block ),
	.I1(\top/processor/seen_last ),
	.I2(\top/processor/n9790_11 ),
	.I3(\top/processor/n11364_28 ),
	.F(\top/processor/n11364_27 )
);
defparam \top/processor/n11364_s21 .INIT=16'h00BF;
LUT4 \top/processor/n11362_s10  (
	.I0(\top/processor/n11362_18 ),
	.I1(\top/processor/n9790_11 ),
	.I2(\top/processor/seen_last ),
	.I3(\top/state_0 [2]),
	.F(\top/processor/n11362_17 )
);
defparam \top/processor/n11362_s10 .INIT=16'hFF40;
LUT4 \top/processor/state_1_s4  (
	.I0(\top/processor/state_1_9 ),
	.I1(\top/processor/n11362_18 ),
	.I2(\top/state_0 [2]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/state_0_10 )
);
defparam \top/processor/state_1_s4 .INIT=16'h030A;
LUT4 \top/processor/byte_index_5_s4  (
	.I0(\top/processor/n8408_6 ),
	.I1(\top/processor/seen_last ),
	.I2(\top/processor/n9790_15 ),
	.I3(\top/processor/total_bits_63_8 ),
	.F(\top/processor/byte_index_5_8 )
);
defparam \top/processor/byte_index_5_s4 .INIT=16'hFF10;
LUT3 \top/processor/core_start_s3  (
	.I0(\top/state_0 [0]),
	.I1(\top/state_0 [1]),
	.I2(\top/state_0 [2]),
	.F(\top/processor/core_start_8 )
);
defparam \top/processor/core_start_s3 .INIT=8'h18;
LUT4 \top/processor/hash_state_255_s4  (
	.I0(\top/processor/n8408_6 ),
	.I1(\top/processor/n9790_11 ),
	.I2(\top/processor/hash_state_255_8 ),
	.I3(\top/state_0 [2]),
	.F(\top/processor/hash_state_255_7 )
);
defparam \top/processor/hash_state_255_s4 .INIT=16'h00F4;
LUT3 \top/processor/total_bits_63_s4  (
	.I0(\top/processor/hash_state_255_8 ),
	.I1(\top/processor/n7631_8 ),
	.I2(\top/state_0 [2]),
	.F(\top/processor/total_bits_63_8 )
);
defparam \top/processor/total_bits_63_s4 .INIT=8'h0E;
LUT4 \top/processor/seen_last_s4  (
	.I0(\top/processor/seen_last_9 ),
	.I1(\top/state_0 [1]),
	.I2(\top/state_0 [2]),
	.I3(\top/data_last ),
	.F(\top/processor/seen_last_8 )
);
defparam \top/processor/seen_last_s4 .INIT=16'h0100;
LUT4 \top/processor/need_length_block_s4  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/need_length_block_9 ),
	.I2(\top/processor/need_length_block_10 ),
	.I3(\top/state_0 [2]),
	.F(\top/processor/need_length_block_8 )
);
defparam \top/processor/need_length_block_s4 .INIT=16'h004F;
LUT4 \top/processor/pad_index_5_s4  (
	.I0(\top/data_last ),
	.I1(\top/state_0 [1]),
	.I2(\top/state_0 [2]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/pad_index_5_8 )
);
defparam \top/processor/pad_index_5_s4 .INIT=16'h000E;
LUT4 \top/processor/block_buffer_503_s4  (
	.I0(\top/processor/block_buffer_503_9 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_503_11 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_503_8 )
);
defparam \top/processor/block_buffer_503_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_495_s4  (
	.I0(\top/processor/block_buffer_495_9 ),
	.I1(\top/processor/block_buffer_495_13 ),
	.I2(\top/processor/block_buffer_495_11 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_495_8 )
);
defparam \top/processor/block_buffer_495_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_487_s4  (
	.I0(\top/processor/block_buffer_495_13 ),
	.I1(\top/processor/block_buffer_487_9 ),
	.I2(\top/processor/block_buffer_487_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_487_8 )
);
defparam \top/processor/block_buffer_487_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_479_s4  (
	.I0(\top/processor/block_buffer_503_9 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_479_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_479_8 )
);
defparam \top/processor/block_buffer_479_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_471_s4  (
	.I0(\top/processor/block_buffer_495_13 ),
	.I1(\top/processor/block_buffer_471_9 ),
	.I2(\top/processor/block_buffer_471_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_471_8 )
);
defparam \top/processor/block_buffer_471_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_463_s4  (
	.I0(\top/processor/block_buffer_495_13 ),
	.I1(\top/processor/block_buffer_463_9 ),
	.I2(\top/processor/block_buffer_463_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_463_8 )
);
defparam \top/processor/block_buffer_463_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_455_s4  (
	.I0(\top/processor/block_buffer_495_13 ),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_455_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_455_8 )
);
defparam \top/processor/block_buffer_455_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_439_s4  (
	.I0(\top/processor/block_buffer_439_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_439_11 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_439_8 )
);
defparam \top/processor/block_buffer_439_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_431_s4  (
	.I0(\top/processor/block_buffer_431_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_431_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_431_8 )
);
defparam \top/processor/block_buffer_431_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_423_s4  (
	.I0(\top/processor/block_buffer_423_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_423_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_423_8 )
);
defparam \top/processor/block_buffer_423_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_415_s4  (
	.I0(\top/processor/block_buffer_415_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_415_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_415_8 )
);
defparam \top/processor/block_buffer_415_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_407_s4  (
	.I0(\top/processor/block_buffer_407_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_407_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_407_8 )
);
defparam \top/processor/block_buffer_407_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_399_s4  (
	.I0(\top/processor/block_buffer_399_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_399_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_399_8 )
);
defparam \top/processor/block_buffer_399_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_391_s4  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/block_buffer_439_10 ),
	.I2(\top/processor/block_buffer_391_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_391_8 )
);
defparam \top/processor/block_buffer_391_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_375_s4  (
	.I0(\top/processor/block_buffer_439_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_375_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_375_8 )
);
defparam \top/processor/block_buffer_375_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_367_s4  (
	.I0(\top/processor/block_buffer_431_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_367_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_367_8 )
);
defparam \top/processor/block_buffer_367_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_359_s4  (
	.I0(\top/processor/block_buffer_423_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_359_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_359_8 )
);
defparam \top/processor/block_buffer_359_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_351_s4  (
	.I0(\top/processor/block_buffer_415_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_351_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_351_8 )
);
defparam \top/processor/block_buffer_351_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_343_s4  (
	.I0(\top/processor/block_buffer_407_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_343_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_343_8 )
);
defparam \top/processor/block_buffer_343_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_335_s4  (
	.I0(\top/processor/block_buffer_399_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_335_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_335_8 )
);
defparam \top/processor/block_buffer_335_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_327_s4  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/block_buffer_375_9 ),
	.I2(\top/processor/block_buffer_327_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_327_8 )
);
defparam \top/processor/block_buffer_327_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_319_s4  (
	.I0(\top/processor/block_buffer_319_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_319_11 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_319_8 )
);
defparam \top/processor/block_buffer_319_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_311_s4  (
	.I0(\top/processor/block_buffer_439_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_311_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_311_8 )
);
defparam \top/processor/block_buffer_311_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_303_s4  (
	.I0(\top/processor/block_buffer_431_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_303_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_303_8 )
);
defparam \top/processor/block_buffer_303_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_295_s4  (
	.I0(\top/processor/block_buffer_423_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_295_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_295_8 )
);
defparam \top/processor/block_buffer_295_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_287_s4  (
	.I0(\top/processor/block_buffer_415_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_287_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_287_8 )
);
defparam \top/processor/block_buffer_287_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_279_s4  (
	.I0(\top/processor/block_buffer_407_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_279_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_279_8 )
);
defparam \top/processor/block_buffer_279_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_271_s4  (
	.I0(\top/processor/block_buffer_399_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_271_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_271_8 )
);
defparam \top/processor/block_buffer_271_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_263_s4  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/block_buffer_319_10 ),
	.I2(\top/processor/block_buffer_263_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_263_8 )
);
defparam \top/processor/block_buffer_263_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_247_s4  (
	.I0(\top/processor/block_buffer_439_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_247_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_247_8 )
);
defparam \top/processor/block_buffer_247_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_239_s4  (
	.I0(\top/processor/block_buffer_431_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_239_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_239_8 )
);
defparam \top/processor/block_buffer_239_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_231_s4  (
	.I0(\top/processor/block_buffer_423_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_231_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_231_8 )
);
defparam \top/processor/block_buffer_231_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_223_s4  (
	.I0(\top/processor/block_buffer_415_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_223_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_223_8 )
);
defparam \top/processor/block_buffer_223_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_215_s4  (
	.I0(\top/processor/block_buffer_407_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_215_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_215_8 )
);
defparam \top/processor/block_buffer_215_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_207_s4  (
	.I0(\top/processor/block_buffer_399_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_207_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_207_8 )
);
defparam \top/processor/block_buffer_207_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_199_s4  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/block_buffer_247_9 ),
	.I2(\top/processor/block_buffer_199_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_199_8 )
);
defparam \top/processor/block_buffer_199_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_191_s4  (
	.I0(\top/processor/block_buffer_319_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_191_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_191_8 )
);
defparam \top/processor/block_buffer_191_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_183_s4  (
	.I0(\top/processor/block_buffer_439_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_183_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_183_8 )
);
defparam \top/processor/block_buffer_183_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_175_s4  (
	.I0(\top/processor/block_buffer_431_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_175_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_175_8 )
);
defparam \top/processor/block_buffer_175_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_167_s4  (
	.I0(\top/processor/block_buffer_423_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_167_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_167_8 )
);
defparam \top/processor/block_buffer_167_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_159_s4  (
	.I0(\top/processor/block_buffer_415_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_159_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_159_8 )
);
defparam \top/processor/block_buffer_159_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_151_s4  (
	.I0(\top/processor/block_buffer_407_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_151_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_151_8 )
);
defparam \top/processor/block_buffer_151_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_143_s4  (
	.I0(\top/processor/block_buffer_399_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_143_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_143_8 )
);
defparam \top/processor/block_buffer_143_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_135_s4  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/block_buffer_191_9 ),
	.I2(\top/processor/block_buffer_135_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_135_8 )
);
defparam \top/processor/block_buffer_135_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_127_s4  (
	.I0(\top/processor/block_buffer_319_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_127_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_127_8 )
);
defparam \top/processor/block_buffer_127_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_119_s4  (
	.I0(\top/processor/block_buffer_439_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_119_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_119_8 )
);
defparam \top/processor/block_buffer_119_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_111_s4  (
	.I0(\top/processor/block_buffer_431_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_111_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_111_8 )
);
defparam \top/processor/block_buffer_111_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_103_s4  (
	.I0(\top/processor/block_buffer_423_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_103_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_103_8 )
);
defparam \top/processor/block_buffer_103_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_95_s4  (
	.I0(\top/processor/block_buffer_415_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_95_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_95_8 )
);
defparam \top/processor/block_buffer_95_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_87_s4  (
	.I0(\top/processor/block_buffer_407_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_87_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_87_8 )
);
defparam \top/processor/block_buffer_87_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_79_s4  (
	.I0(\top/processor/block_buffer_399_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_79_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_79_8 )
);
defparam \top/processor/block_buffer_79_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_71_s4  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/block_buffer_127_9 ),
	.I2(\top/processor/block_buffer_71_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_71_8 )
);
defparam \top/processor/block_buffer_71_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_63_s4  (
	.I0(\top/processor/block_buffer_63_9 ),
	.I1(\top/processor/block_buffer_63_10 ),
	.I2(\top/processor/block_buffer_63_11 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_63_8 )
);
defparam \top/processor/block_buffer_63_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_55_s4  (
	.I0(\top/processor/block_buffer_55_9 ),
	.I1(\top/processor/block_buffer_55_10 ),
	.I2(\top/processor/n7631_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_55_8 )
);
defparam \top/processor/block_buffer_55_s4 .INIT=16'hEF00;
LUT4 \top/processor/block_buffer_47_s4  (
	.I0(\top/processor/block_buffer_63_9 ),
	.I1(\top/processor/block_buffer_495_9 ),
	.I2(\top/processor/block_buffer_47_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_47_8 )
);
defparam \top/processor/block_buffer_47_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_39_s4  (
	.I0(\top/processor/block_buffer_63_9 ),
	.I1(\top/processor/block_buffer_487_9 ),
	.I2(\top/processor/block_buffer_39_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_39_8 )
);
defparam \top/processor/block_buffer_39_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_31_s4  (
	.I0(\top/processor/block_buffer_31_9 ),
	.I1(\top/processor/block_buffer_31_10 ),
	.I2(\top/processor/n7631_10 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_31_8 )
);
defparam \top/processor/block_buffer_31_s4 .INIT=16'hEF00;
LUT4 \top/processor/block_buffer_23_s4  (
	.I0(\top/processor/block_buffer_63_9 ),
	.I1(\top/processor/block_buffer_471_9 ),
	.I2(\top/processor/block_buffer_23_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_23_8 )
);
defparam \top/processor/block_buffer_23_s4 .INIT=16'h8F00;
LUT4 \top/processor/block_buffer_15_s4  (
	.I0(\top/processor/block_buffer_63_9 ),
	.I1(\top/processor/block_buffer_463_9 ),
	.I2(\top/processor/block_buffer_15_9 ),
	.I3(\top/processor/block_buffer_511_11 ),
	.F(\top/processor/block_buffer_15_8 )
);
defparam \top/processor/block_buffer_15_s4 .INIT=16'h8F00;
LUT3 \top/processor/block_ready_s4  (
	.I0(\top/state_0 [2]),
	.I1(\top/processor/n7631_3 ),
	.I2(\top/processor/n9790_13 ),
	.F(\top/processor/block_ready_8 )
);
defparam \top/processor/block_ready_s4 .INIT=8'hF4;
LUT2 \top/processor/n11438_s9  (
	.I0(\top/processor/total_bits [3]),
	.I1(\top/state_0 [0]),
	.F(\top/processor/n11438_14 )
);
defparam \top/processor/n11438_s9 .INIT=4'h4;
LUT3 \top/processor/n11437_s9  (
	.I0(\top/processor/total_bits [4]),
	.I1(\top/processor/total_bits [3]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11437_14 )
);
defparam \top/processor/n11437_s9 .INIT=8'h60;
LUT4 \top/processor/n11436_s9  (
	.I0(\top/processor/total_bits [4]),
	.I1(\top/processor/total_bits [3]),
	.I2(\top/processor/total_bits [5]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11436_14 )
);
defparam \top/processor/n11436_s9 .INIT=16'h7800;
LUT3 \top/processor/n11435_s9  (
	.I0(\top/processor/n11435_15 ),
	.I1(\top/processor/total_bits [6]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11435_14 )
);
defparam \top/processor/n11435_s9 .INIT=8'h60;
LUT3 \top/processor/n11434_s9  (
	.I0(\top/processor/total_bits [7]),
	.I1(\top/processor/n11434_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11434_14 )
);
defparam \top/processor/n11434_s9 .INIT=8'h60;
LUT4 \top/processor/n11433_s9  (
	.I0(\top/processor/total_bits [7]),
	.I1(\top/processor/n11434_15 ),
	.I2(\top/processor/total_bits [8]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11433_14 )
);
defparam \top/processor/n11433_s9 .INIT=16'h7800;
LUT3 \top/processor/n11432_s9  (
	.I0(\top/processor/n11432_15 ),
	.I1(\top/processor/total_bits [9]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11432_14 )
);
defparam \top/processor/n11432_s9 .INIT=8'h60;
LUT3 \top/processor/n11431_s9  (
	.I0(\top/processor/total_bits [10]),
	.I1(\top/processor/n11431_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11431_14 )
);
defparam \top/processor/n11431_s9 .INIT=8'h60;
LUT4 \top/processor/n11429_s9  (
	.I0(\top/processor/total_bits [11]),
	.I1(\top/processor/n11430_15 ),
	.I2(\top/processor/total_bits [12]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11429_14 )
);
defparam \top/processor/n11429_s9 .INIT=16'h7800;
LUT4 \top/processor/n11428_s9  (
	.I0(\top/processor/n11430_15 ),
	.I1(\top/processor/n11428_15 ),
	.I2(\top/processor/total_bits [13]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11428_14 )
);
defparam \top/processor/n11428_s9 .INIT=16'h7800;
LUT3 \top/processor/n11427_s9  (
	.I0(\top/processor/total_bits [14]),
	.I1(\top/processor/n11427_17 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11427_14 )
);
defparam \top/processor/n11427_s9 .INIT=8'h60;
LUT4 \top/processor/n11426_s9  (
	.I0(\top/processor/total_bits [14]),
	.I1(\top/processor/n11427_17 ),
	.I2(\top/processor/total_bits [15]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11426_14 )
);
defparam \top/processor/n11426_s9 .INIT=16'h7800;
LUT4 \top/processor/n11425_s9  (
	.I0(\top/processor/n11430_15 ),
	.I1(\top/processor/n11425_15 ),
	.I2(\top/processor/total_bits [16]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11425_14 )
);
defparam \top/processor/n11425_s9 .INIT=16'h7800;
LUT3 \top/processor/n11424_s9  (
	.I0(\top/processor/total_bits [17]),
	.I1(\top/processor/n11424_17 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11424_14 )
);
defparam \top/processor/n11424_s9 .INIT=8'h60;
LUT4 \top/processor/n11422_s9  (
	.I0(\top/processor/total_bits [18]),
	.I1(\top/processor/n11423_15 ),
	.I2(\top/processor/total_bits [19]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11422_14 )
);
defparam \top/processor/n11422_s9 .INIT=16'h7800;
LUT3 \top/processor/n11421_s9  (
	.I0(\top/processor/n11421_17 ),
	.I1(\top/processor/total_bits [20]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11421_14 )
);
defparam \top/processor/n11421_s9 .INIT=8'h60;
LUT3 \top/processor/n11420_s9  (
	.I0(\top/processor/total_bits [21]),
	.I1(\top/processor/n11420_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11420_14 )
);
defparam \top/processor/n11420_s9 .INIT=8'h60;
LUT4 \top/processor/n11419_s9  (
	.I0(\top/processor/total_bits [21]),
	.I1(\top/processor/n11420_15 ),
	.I2(\top/processor/total_bits [22]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11419_14 )
);
defparam \top/processor/n11419_s9 .INIT=16'h7800;
LUT3 \top/processor/n11418_s9  (
	.I0(\top/processor/n11418_15 ),
	.I1(\top/processor/total_bits [23]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11418_14 )
);
defparam \top/processor/n11418_s9 .INIT=8'h60;
LUT4 \top/processor/n11417_s9  (
	.I0(\top/processor/n11420_15 ),
	.I1(\top/processor/n11417_15 ),
	.I2(\top/processor/total_bits [24]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11417_14 )
);
defparam \top/processor/n11417_s9 .INIT=16'h7800;
LUT3 \top/processor/n11416_s9  (
	.I0(\top/processor/n11416_15 ),
	.I1(\top/processor/total_bits [25]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11416_14 )
);
defparam \top/processor/n11416_s9 .INIT=8'h60;
LUT3 \top/processor/n11415_s9  (
	.I0(\top/processor/total_bits [26]),
	.I1(\top/processor/n11415_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11415_14 )
);
defparam \top/processor/n11415_s9 .INIT=8'h60;
LUT4 \top/processor/n11413_s9  (
	.I0(\top/processor/total_bits [27]),
	.I1(\top/processor/n11414_15 ),
	.I2(\top/processor/total_bits [28]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11413_14 )
);
defparam \top/processor/n11413_s9 .INIT=16'h7800;
LUT4 \top/processor/n11412_s9  (
	.I0(\top/processor/n11414_15 ),
	.I1(\top/processor/n11412_15 ),
	.I2(\top/processor/total_bits [29]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11412_14 )
);
defparam \top/processor/n11412_s9 .INIT=16'h7800;
LUT4 \top/processor/n11411_s9  (
	.I0(\top/processor/n11414_15 ),
	.I1(\top/processor/n11411_15 ),
	.I2(\top/processor/total_bits [30]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11411_14 )
);
defparam \top/processor/n11411_s9 .INIT=16'h7800;
LUT3 \top/processor/n11410_s9  (
	.I0(\top/processor/total_bits [31]),
	.I1(\top/processor/n11410_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11410_14 )
);
defparam \top/processor/n11410_s9 .INIT=8'h60;
LUT4 \top/processor/n11408_s9  (
	.I0(\top/processor/total_bits [32]),
	.I1(\top/processor/n11409_15 ),
	.I2(\top/processor/total_bits [33]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11408_14 )
);
defparam \top/processor/n11408_s9 .INIT=16'h7800;
LUT3 \top/processor/n11407_s9  (
	.I0(\top/processor/total_bits [34]),
	.I1(\top/processor/n11407_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11407_14 )
);
defparam \top/processor/n11407_s9 .INIT=8'h60;
LUT4 \top/processor/n11406_s9  (
	.I0(\top/processor/total_bits [34]),
	.I1(\top/processor/n11407_15 ),
	.I2(\top/processor/total_bits [35]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11406_14 )
);
defparam \top/processor/n11406_s9 .INIT=16'h7800;
LUT3 \top/processor/n11405_s9  (
	.I0(\top/processor/total_bits [36]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11405_14 )
);
defparam \top/processor/n11405_s9 .INIT=8'h60;
LUT4 \top/processor/n11404_s9  (
	.I0(\top/processor/total_bits [36]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/total_bits [37]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11404_14 )
);
defparam \top/processor/n11404_s9 .INIT=16'h7800;
LUT4 \top/processor/n11403_s9  (
	.I0(\top/processor/n11405_15 ),
	.I1(\top/processor/n11403_15 ),
	.I2(\top/processor/total_bits [38]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11403_14 )
);
defparam \top/processor/n11403_s9 .INIT=16'h7800;
LUT3 \top/processor/n11402_s9  (
	.I0(\top/processor/total_bits [39]),
	.I1(\top/processor/n11402_17 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11402_14 )
);
defparam \top/processor/n11402_s9 .INIT=8'h60;
LUT4 \top/processor/n11401_s9  (
	.I0(\top/processor/total_bits [39]),
	.I1(\top/processor/n11402_17 ),
	.I2(\top/processor/total_bits [40]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11401_14 )
);
defparam \top/processor/n11401_s9 .INIT=16'h7800;
LUT4 \top/processor/n11400_s9  (
	.I0(\top/processor/n11405_15 ),
	.I1(\top/processor/n11400_15 ),
	.I2(\top/processor/total_bits [41]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11400_14 )
);
defparam \top/processor/n11400_s9 .INIT=16'h7800;
LUT3 \top/processor/n11399_s9  (
	.I0(\top/processor/n11399_15 ),
	.I1(\top/processor/total_bits [42]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11399_14 )
);
defparam \top/processor/n11399_s9 .INIT=8'h60;
LUT3 \top/processor/n11398_s9  (
	.I0(\top/processor/total_bits [43]),
	.I1(\top/processor/n11398_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11398_14 )
);
defparam \top/processor/n11398_s9 .INIT=8'h60;
LUT4 \top/processor/n11397_s9  (
	.I0(\top/processor/total_bits [43]),
	.I1(\top/processor/n11398_15 ),
	.I2(\top/processor/total_bits [44]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11397_14 )
);
defparam \top/processor/n11397_s9 .INIT=16'h7800;
LUT3 \top/processor/n11396_s9  (
	.I0(\top/processor/n11396_15 ),
	.I1(\top/processor/total_bits [45]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11396_14 )
);
defparam \top/processor/n11396_s9 .INIT=8'h60;
LUT4 \top/processor/n11395_s9  (
	.I0(\top/processor/n11405_15 ),
	.I1(\top/processor/n11395_15 ),
	.I2(\top/processor/total_bits [46]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11395_14 )
);
defparam \top/processor/n11395_s9 .INIT=16'h7800;
LUT3 \top/processor/n11394_s9  (
	.I0(\top/processor/total_bits [47]),
	.I1(\top/processor/n11394_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11394_14 )
);
defparam \top/processor/n11394_s9 .INIT=8'h60;
LUT4 \top/processor/n11393_s9  (
	.I0(\top/processor/total_bits [47]),
	.I1(\top/processor/n11394_15 ),
	.I2(\top/processor/total_bits [48]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11393_14 )
);
defparam \top/processor/n11393_s9 .INIT=16'h7800;
LUT3 \top/processor/n11392_s9  (
	.I0(\top/processor/total_bits [49]),
	.I1(\top/processor/n11392_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11392_14 )
);
defparam \top/processor/n11392_s9 .INIT=8'h60;
LUT4 \top/processor/n11391_s9  (
	.I0(\top/processor/total_bits [49]),
	.I1(\top/processor/n11392_15 ),
	.I2(\top/processor/total_bits [50]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11391_14 )
);
defparam \top/processor/n11391_s9 .INIT=16'h7800;
LUT4 \top/processor/n11389_s9  (
	.I0(\top/processor/total_bits [51]),
	.I1(\top/processor/n11390_15 ),
	.I2(\top/processor/total_bits [52]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11389_14 )
);
defparam \top/processor/n11389_s9 .INIT=16'h7800;
LUT4 \top/processor/n11388_s9  (
	.I0(\top/processor/n11390_15 ),
	.I1(\top/processor/n11388_15 ),
	.I2(\top/processor/total_bits [53]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11388_14 )
);
defparam \top/processor/n11388_s9 .INIT=16'h7800;
LUT3 \top/processor/n11387_s9  (
	.I0(\top/processor/total_bits [54]),
	.I1(\top/processor/n11387_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11387_14 )
);
defparam \top/processor/n11387_s9 .INIT=8'h60;
LUT4 \top/processor/n11386_s9  (
	.I0(\top/processor/total_bits [54]),
	.I1(\top/processor/n11387_15 ),
	.I2(\top/processor/total_bits [55]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11386_14 )
);
defparam \top/processor/n11386_s9 .INIT=16'h7800;
LUT3 \top/processor/n11385_s9  (
	.I0(\top/processor/total_bits [56]),
	.I1(\top/processor/n11385_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11385_14 )
);
defparam \top/processor/n11385_s9 .INIT=8'h60;
LUT4 \top/processor/n11384_s9  (
	.I0(\top/processor/total_bits [56]),
	.I1(\top/processor/n11385_15 ),
	.I2(\top/processor/total_bits [57]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11384_14 )
);
defparam \top/processor/n11384_s9 .INIT=16'h7800;
LUT4 \top/processor/n11383_s9  (
	.I0(\top/processor/n11385_15 ),
	.I1(\top/processor/n11383_15 ),
	.I2(\top/processor/total_bits [58]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11383_14 )
);
defparam \top/processor/n11383_s9 .INIT=16'h7800;
LUT3 \top/processor/n11382_s9  (
	.I0(\top/processor/total_bits [59]),
	.I1(\top/processor/n11382_15 ),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11382_14 )
);
defparam \top/processor/n11382_s9 .INIT=8'h60;
LUT4 \top/processor/n11381_s9  (
	.I0(\top/processor/total_bits [59]),
	.I1(\top/processor/n11382_15 ),
	.I2(\top/processor/total_bits [60]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11381_14 )
);
defparam \top/processor/n11381_s9 .INIT=16'h7800;
LUT4 \top/processor/n11380_s9  (
	.I0(\top/processor/n11382_15 ),
	.I1(\top/processor/n11380_15 ),
	.I2(\top/processor/total_bits [61]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11380_14 )
);
defparam \top/processor/n11380_s9 .INIT=16'h7800;
LUT4 \top/processor/n11379_s9  (
	.I0(\top/processor/n11382_15 ),
	.I1(\top/processor/n11379_17 ),
	.I2(\top/processor/total_bits [62]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11379_14 )
);
defparam \top/processor/n11379_s9 .INIT=16'h7800;
LUT4 \top/processor/n11378_s9  (
	.I0(\top/processor/n11382_15 ),
	.I1(\top/processor/n11378_17 ),
	.I2(\top/processor/total_bits [63]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11378_14 )
);
defparam \top/processor/n11378_s9 .INIT=16'h7800;
LUT4 \top/processor/n11377_s9  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/n11377_15 ),
	.I2(\top/processor/n10817_15 ),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11377_14 )
);
defparam \top/processor/n11377_s9 .INIT=16'h5C00;
LUT2 \top/processor/n11376_s9  (
	.I0(\top/processor/n11376_15 ),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n11376_14 )
);
defparam \top/processor/n11376_s9 .INIT=4'h4;
LUT4 \top/processor/n11375_s9  (
	.I0(\top/processor/n11375_15 ),
	.I1(\top/processor/n10817_15 ),
	.I2(\top/processor/n11375_16 ),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11375_14 )
);
defparam \top/processor/n11375_s9 .INIT=16'hF800;
LUT4 \top/processor/n11374_s9  (
	.I0(\top/processor/n11374_20 ),
	.I1(\top/processor/n11374_22 ),
	.I2(\top/processor/n11374_17 ),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11374_14 )
);
defparam \top/processor/n11374_s9 .INIT=16'hF400;
LUT4 \top/processor/n11373_s9  (
	.I0(\top/processor/n11373_15 ),
	.I1(\top/processor/n10817_15 ),
	.I2(\top/processor/n11373_16 ),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11373_14 )
);
defparam \top/processor/n11373_s9 .INIT=16'hF800;
LUT4 \top/processor/n11372_s9  (
	.I0(\top/processor/n10817_15 ),
	.I1(\top/processor/n11372_15 ),
	.I2(\top/processor/n11372_16 ),
	.I3(\top/state_0 [1]),
	.F(\top/processor/n11372_14 )
);
defparam \top/processor/n11372_s9 .INIT=16'h2F00;
LUT4 \top/processor/n11368_s11  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [2]),
	.I3(\top/processor/n11370_19 ),
	.F(\top/processor/n11368_17 )
);
defparam \top/processor/n11368_s11 .INIT=16'h7800;
LUT4 \top/processor/n11366_s11  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/block_buffer_391_9 ),
	.I2(\top/processor/byte_index [4]),
	.I3(\top/processor/n11370_19 ),
	.F(\top/processor/n11366_17 )
);
defparam \top/processor/n11366_s11 .INIT=16'h7800;
LUT2 \top/processor/n10824_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [0]),
	.F(\top/processor/n10824_15 )
);
defparam \top/processor/n10824_s10 .INIT=4'h4;
LUT2 \top/processor/n10823_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [1]),
	.F(\top/processor/n10823_15 )
);
defparam \top/processor/n10823_s10 .INIT=4'h4;
LUT2 \top/processor/n10822_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [2]),
	.F(\top/processor/n10822_15 )
);
defparam \top/processor/n10822_s10 .INIT=4'h4;
LUT2 \top/processor/n10821_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [3]),
	.F(\top/processor/n10821_15 )
);
defparam \top/processor/n10821_s10 .INIT=4'h4;
LUT2 \top/processor/n10820_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [4]),
	.F(\top/processor/n10820_15 )
);
defparam \top/processor/n10820_s10 .INIT=4'h4;
LUT2 \top/processor/n10819_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [5]),
	.F(\top/processor/n10819_15 )
);
defparam \top/processor/n10819_s10 .INIT=4'h4;
LUT2 \top/processor/n10818_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/data_in [6]),
	.F(\top/processor/n10818_15 )
);
defparam \top/processor/n10818_s10 .INIT=4'h4;
LUT2 \top/processor/n10815_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [1]),
	.F(\top/processor/n10815_15 )
);
defparam \top/processor/n10815_s10 .INIT=4'h8;
LUT2 \top/processor/n10814_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [2]),
	.F(\top/processor/n10814_15 )
);
defparam \top/processor/n10814_s10 .INIT=4'h8;
LUT2 \top/processor/n10811_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [5]),
	.F(\top/processor/n10811_15 )
);
defparam \top/processor/n10811_s10 .INIT=4'h8;
LUT2 \top/processor/n10810_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [6]),
	.F(\top/processor/n10810_15 )
);
defparam \top/processor/n10810_s10 .INIT=4'h8;
LUT2 \top/processor/n10809_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [7]),
	.F(\top/processor/n10809_15 )
);
defparam \top/processor/n10809_s10 .INIT=4'h8;
LUT2 \top/processor/n10807_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [9]),
	.F(\top/processor/n10807_15 )
);
defparam \top/processor/n10807_s10 .INIT=4'h8;
LUT2 \top/processor/n10804_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [12]),
	.F(\top/processor/n10804_15 )
);
defparam \top/processor/n10804_s10 .INIT=4'h8;
LUT2 \top/processor/n10803_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [13]),
	.F(\top/processor/n10803_15 )
);
defparam \top/processor/n10803_s10 .INIT=4'h8;
LUT2 \top/processor/n10800_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [16]),
	.F(\top/processor/n10800_15 )
);
defparam \top/processor/n10800_s10 .INIT=4'h8;
LUT2 \top/processor/n10799_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [17]),
	.F(\top/processor/n10799_15 )
);
defparam \top/processor/n10799_s10 .INIT=4'h8;
LUT2 \top/processor/n10798_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [18]),
	.F(\top/processor/n10798_15 )
);
defparam \top/processor/n10798_s10 .INIT=4'h8;
LUT2 \top/processor/n10797_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [19]),
	.F(\top/processor/n10797_15 )
);
defparam \top/processor/n10797_s10 .INIT=4'h8;
LUT2 \top/processor/n10796_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [20]),
	.F(\top/processor/n10796_15 )
);
defparam \top/processor/n10796_s10 .INIT=4'h8;
LUT2 \top/processor/n10790_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [26]),
	.F(\top/processor/n10790_15 )
);
defparam \top/processor/n10790_s10 .INIT=4'h8;
LUT2 \top/processor/n10787_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [29]),
	.F(\top/processor/n10787_15 )
);
defparam \top/processor/n10787_s10 .INIT=4'h8;
LUT2 \top/processor/n10785_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [31]),
	.F(\top/processor/n10785_15 )
);
defparam \top/processor/n10785_s10 .INIT=4'h8;
LUT2 \top/processor/n10782_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [34]),
	.F(\top/processor/n10782_15 )
);
defparam \top/processor/n10782_s10 .INIT=4'h8;
LUT2 \top/processor/n10780_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [36]),
	.F(\top/processor/n10780_15 )
);
defparam \top/processor/n10780_s10 .INIT=4'h8;
LUT2 \top/processor/n10778_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [38]),
	.F(\top/processor/n10778_15 )
);
defparam \top/processor/n10778_s10 .INIT=4'h8;
LUT2 \top/processor/n10775_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [41]),
	.F(\top/processor/n10775_15 )
);
defparam \top/processor/n10775_s10 .INIT=4'h8;
LUT2 \top/processor/n10774_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [42]),
	.F(\top/processor/n10774_15 )
);
defparam \top/processor/n10774_s10 .INIT=4'h8;
LUT2 \top/processor/n10771_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [45]),
	.F(\top/processor/n10771_15 )
);
defparam \top/processor/n10771_s10 .INIT=4'h8;
LUT2 \top/processor/n10766_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [50]),
	.F(\top/processor/n10766_15 )
);
defparam \top/processor/n10766_s10 .INIT=4'h8;
LUT2 \top/processor/n10765_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [51]),
	.F(\top/processor/n10765_15 )
);
defparam \top/processor/n10765_s10 .INIT=4'h8;
LUT2 \top/processor/n10764_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [52]),
	.F(\top/processor/n10764_15 )
);
defparam \top/processor/n10764_s10 .INIT=4'h8;
LUT2 \top/processor/n10763_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [53]),
	.F(\top/processor/n10763_15 )
);
defparam \top/processor/n10763_s10 .INIT=4'h8;
LUT2 \top/processor/n10762_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [54]),
	.F(\top/processor/n10762_15 )
);
defparam \top/processor/n10762_s10 .INIT=4'h8;
LUT2 \top/processor/n10755_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [61]),
	.F(\top/processor/n10755_15 )
);
defparam \top/processor/n10755_s10 .INIT=4'h8;
LUT2 \top/processor/n10754_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [62]),
	.F(\top/processor/n10754_15 )
);
defparam \top/processor/n10754_s10 .INIT=4'h8;
LUT2 \top/processor/n10753_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [63]),
	.F(\top/processor/n10753_15 )
);
defparam \top/processor/n10753_s10 .INIT=4'h8;
LUT2 \top/processor/n10752_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [64]),
	.F(\top/processor/n10752_15 )
);
defparam \top/processor/n10752_s10 .INIT=4'h8;
LUT2 \top/processor/n10751_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [65]),
	.F(\top/processor/n10751_15 )
);
defparam \top/processor/n10751_s10 .INIT=4'h8;
LUT2 \top/processor/n10748_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [68]),
	.F(\top/processor/n10748_15 )
);
defparam \top/processor/n10748_s10 .INIT=4'h8;
LUT2 \top/processor/n10747_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [69]),
	.F(\top/processor/n10747_15 )
);
defparam \top/processor/n10747_s10 .INIT=4'h8;
LUT2 \top/processor/n10746_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [70]),
	.F(\top/processor/n10746_15 )
);
defparam \top/processor/n10746_s10 .INIT=4'h8;
LUT2 \top/processor/n10744_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [72]),
	.F(\top/processor/n10744_15 )
);
defparam \top/processor/n10744_s10 .INIT=4'h8;
LUT2 \top/processor/n10743_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [73]),
	.F(\top/processor/n10743_15 )
);
defparam \top/processor/n10743_s10 .INIT=4'h8;
LUT2 \top/processor/n10742_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [74]),
	.F(\top/processor/n10742_15 )
);
defparam \top/processor/n10742_s10 .INIT=4'h8;
LUT2 \top/processor/n10740_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [76]),
	.F(\top/processor/n10740_15 )
);
defparam \top/processor/n10740_s10 .INIT=4'h8;
LUT2 \top/processor/n10737_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [79]),
	.F(\top/processor/n10737_15 )
);
defparam \top/processor/n10737_s10 .INIT=4'h8;
LUT2 \top/processor/n10735_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [81]),
	.F(\top/processor/n10735_15 )
);
defparam \top/processor/n10735_s10 .INIT=4'h8;
LUT2 \top/processor/n10733_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [83]),
	.F(\top/processor/n10733_15 )
);
defparam \top/processor/n10733_s10 .INIT=4'h8;
LUT2 \top/processor/n10732_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [84]),
	.F(\top/processor/n10732_15 )
);
defparam \top/processor/n10732_s10 .INIT=4'h8;
LUT2 \top/processor/n10731_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [85]),
	.F(\top/processor/n10731_15 )
);
defparam \top/processor/n10731_s10 .INIT=4'h8;
LUT2 \top/processor/n10730_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [86]),
	.F(\top/processor/n10730_15 )
);
defparam \top/processor/n10730_s10 .INIT=4'h8;
LUT2 \top/processor/n10729_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [87]),
	.F(\top/processor/n10729_15 )
);
defparam \top/processor/n10729_s10 .INIT=4'h8;
LUT2 \top/processor/n10726_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [90]),
	.F(\top/processor/n10726_15 )
);
defparam \top/processor/n10726_s10 .INIT=4'h8;
LUT2 \top/processor/n10723_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [93]),
	.F(\top/processor/n10723_15 )
);
defparam \top/processor/n10723_s10 .INIT=4'h8;
LUT2 \top/processor/n10722_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [94]),
	.F(\top/processor/n10722_15 )
);
defparam \top/processor/n10722_s10 .INIT=4'h8;
LUT2 \top/processor/n10713_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [103]),
	.F(\top/processor/n10713_15 )
);
defparam \top/processor/n10713_s10 .INIT=4'h8;
LUT2 \top/processor/n10712_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [104]),
	.F(\top/processor/n10712_15 )
);
defparam \top/processor/n10712_s10 .INIT=4'h8;
LUT2 \top/processor/n10710_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [106]),
	.F(\top/processor/n10710_15 )
);
defparam \top/processor/n10710_s10 .INIT=4'h8;
LUT2 \top/processor/n10709_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [107]),
	.F(\top/processor/n10709_15 )
);
defparam \top/processor/n10709_s10 .INIT=4'h8;
LUT2 \top/processor/n10707_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [109]),
	.F(\top/processor/n10707_15 )
);
defparam \top/processor/n10707_s10 .INIT=4'h8;
LUT2 \top/processor/n10705_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [111]),
	.F(\top/processor/n10705_15 )
);
defparam \top/processor/n10705_s10 .INIT=4'h8;
LUT2 \top/processor/n10704_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [112]),
	.F(\top/processor/n10704_15 )
);
defparam \top/processor/n10704_s10 .INIT=4'h8;
LUT2 \top/processor/n10700_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [116]),
	.F(\top/processor/n10700_15 )
);
defparam \top/processor/n10700_s10 .INIT=4'h8;
LUT2 \top/processor/n10699_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [117]),
	.F(\top/processor/n10699_15 )
);
defparam \top/processor/n10699_s10 .INIT=4'h8;
LUT2 \top/processor/n10698_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [118]),
	.F(\top/processor/n10698_15 )
);
defparam \top/processor/n10698_s10 .INIT=4'h8;
LUT2 \top/processor/n10697_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [119]),
	.F(\top/processor/n10697_15 )
);
defparam \top/processor/n10697_s10 .INIT=4'h8;
LUT2 \top/processor/n10695_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [121]),
	.F(\top/processor/n10695_15 )
);
defparam \top/processor/n10695_s10 .INIT=4'h8;
LUT2 \top/processor/n10694_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [122]),
	.F(\top/processor/n10694_15 )
);
defparam \top/processor/n10694_s10 .INIT=4'h8;
LUT2 \top/processor/n10693_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [123]),
	.F(\top/processor/n10693_15 )
);
defparam \top/processor/n10693_s10 .INIT=4'h8;
LUT2 \top/processor/n10691_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [125]),
	.F(\top/processor/n10691_15 )
);
defparam \top/processor/n10691_s10 .INIT=4'h8;
LUT2 \top/processor/n10689_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [127]),
	.F(\top/processor/n10689_15 )
);
defparam \top/processor/n10689_s10 .INIT=4'h8;
LUT2 \top/processor/n10688_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [128]),
	.F(\top/processor/n10688_15 )
);
defparam \top/processor/n10688_s10 .INIT=4'h8;
LUT2 \top/processor/n10686_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [130]),
	.F(\top/processor/n10686_15 )
);
defparam \top/processor/n10686_s10 .INIT=4'h8;
LUT2 \top/processor/n10682_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [134]),
	.F(\top/processor/n10682_15 )
);
defparam \top/processor/n10682_s10 .INIT=4'h8;
LUT2 \top/processor/n10681_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [135]),
	.F(\top/processor/n10681_15 )
);
defparam \top/processor/n10681_s10 .INIT=4'h8;
LUT2 \top/processor/n10679_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [137]),
	.F(\top/processor/n10679_15 )
);
defparam \top/processor/n10679_s10 .INIT=4'h8;
LUT2 \top/processor/n10677_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [139]),
	.F(\top/processor/n10677_15 )
);
defparam \top/processor/n10677_s10 .INIT=4'h8;
LUT2 \top/processor/n10668_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [148]),
	.F(\top/processor/n10668_15 )
);
defparam \top/processor/n10668_s10 .INIT=4'h8;
LUT2 \top/processor/n10667_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [149]),
	.F(\top/processor/n10667_15 )
);
defparam \top/processor/n10667_s10 .INIT=4'h8;
LUT2 \top/processor/n10665_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [151]),
	.F(\top/processor/n10665_15 )
);
defparam \top/processor/n10665_s10 .INIT=4'h8;
LUT2 \top/processor/n10663_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [153]),
	.F(\top/processor/n10663_15 )
);
defparam \top/processor/n10663_s10 .INIT=4'h8;
LUT2 \top/processor/n10661_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [155]),
	.F(\top/processor/n10661_15 )
);
defparam \top/processor/n10661_s10 .INIT=4'h8;
LUT2 \top/processor/n10660_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [156]),
	.F(\top/processor/n10660_15 )
);
defparam \top/processor/n10660_s10 .INIT=4'h8;
LUT2 \top/processor/n10658_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [158]),
	.F(\top/processor/n10658_15 )
);
defparam \top/processor/n10658_s10 .INIT=4'h8;
LUT2 \top/processor/n10656_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [160]),
	.F(\top/processor/n10656_15 )
);
defparam \top/processor/n10656_s10 .INIT=4'h8;
LUT2 \top/processor/n10654_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [162]),
	.F(\top/processor/n10654_15 )
);
defparam \top/processor/n10654_s10 .INIT=4'h8;
LUT2 \top/processor/n10653_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [163]),
	.F(\top/processor/n10653_15 )
);
defparam \top/processor/n10653_s10 .INIT=4'h8;
LUT2 \top/processor/n10649_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [167]),
	.F(\top/processor/n10649_15 )
);
defparam \top/processor/n10649_s10 .INIT=4'h8;
LUT2 \top/processor/n10646_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [170]),
	.F(\top/processor/n10646_15 )
);
defparam \top/processor/n10646_s10 .INIT=4'h8;
LUT2 \top/processor/n10645_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [171]),
	.F(\top/processor/n10645_15 )
);
defparam \top/processor/n10645_s10 .INIT=4'h8;
LUT2 \top/processor/n10640_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [176]),
	.F(\top/processor/n10640_15 )
);
defparam \top/processor/n10640_s10 .INIT=4'h8;
LUT2 \top/processor/n10636_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [180]),
	.F(\top/processor/n10636_15 )
);
defparam \top/processor/n10636_s10 .INIT=4'h8;
LUT2 \top/processor/n10633_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [183]),
	.F(\top/processor/n10633_15 )
);
defparam \top/processor/n10633_s10 .INIT=4'h8;
LUT2 \top/processor/n10632_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [184]),
	.F(\top/processor/n10632_15 )
);
defparam \top/processor/n10632_s10 .INIT=4'h8;
LUT2 \top/processor/n10631_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [185]),
	.F(\top/processor/n10631_15 )
);
defparam \top/processor/n10631_s10 .INIT=4'h8;
LUT2 \top/processor/n10626_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [190]),
	.F(\top/processor/n10626_15 )
);
defparam \top/processor/n10626_s10 .INIT=4'h8;
LUT2 \top/processor/n10625_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [191]),
	.F(\top/processor/n10625_15 )
);
defparam \top/processor/n10625_s10 .INIT=4'h8;
LUT2 \top/processor/n10623_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [193]),
	.F(\top/processor/n10623_15 )
);
defparam \top/processor/n10623_s10 .INIT=4'h8;
LUT2 \top/processor/n10621_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [195]),
	.F(\top/processor/n10621_15 )
);
defparam \top/processor/n10621_s10 .INIT=4'h8;
LUT2 \top/processor/n10620_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [196]),
	.F(\top/processor/n10620_15 )
);
defparam \top/processor/n10620_s10 .INIT=4'h8;
LUT2 \top/processor/n10619_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [197]),
	.F(\top/processor/n10619_15 )
);
defparam \top/processor/n10619_s10 .INIT=4'h8;
LUT2 \top/processor/n10618_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [198]),
	.F(\top/processor/n10618_15 )
);
defparam \top/processor/n10618_s10 .INIT=4'h8;
LUT2 \top/processor/n10616_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [200]),
	.F(\top/processor/n10616_15 )
);
defparam \top/processor/n10616_s10 .INIT=4'h8;
LUT2 \top/processor/n10612_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [204]),
	.F(\top/processor/n10612_15 )
);
defparam \top/processor/n10612_s10 .INIT=4'h8;
LUT2 \top/processor/n10610_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [206]),
	.F(\top/processor/n10610_15 )
);
defparam \top/processor/n10610_s10 .INIT=4'h8;
LUT2 \top/processor/n10605_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [211]),
	.F(\top/processor/n10605_15 )
);
defparam \top/processor/n10605_s10 .INIT=4'h8;
LUT2 \top/processor/n10604_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [212]),
	.F(\top/processor/n10604_15 )
);
defparam \top/processor/n10604_s10 .INIT=4'h8;
LUT2 \top/processor/n10601_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [215]),
	.F(\top/processor/n10601_15 )
);
defparam \top/processor/n10601_s10 .INIT=4'h8;
LUT2 \top/processor/n10598_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [218]),
	.F(\top/processor/n10598_15 )
);
defparam \top/processor/n10598_s10 .INIT=4'h8;
LUT2 \top/processor/n10594_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [222]),
	.F(\top/processor/n10594_15 )
);
defparam \top/processor/n10594_s10 .INIT=4'h8;
LUT2 \top/processor/n10589_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [227]),
	.F(\top/processor/n10589_15 )
);
defparam \top/processor/n10589_s10 .INIT=4'h8;
LUT2 \top/processor/n10588_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [228]),
	.F(\top/processor/n10588_15 )
);
defparam \top/processor/n10588_s10 .INIT=4'h8;
LUT2 \top/processor/n10585_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [231]),
	.F(\top/processor/n10585_15 )
);
defparam \top/processor/n10585_s10 .INIT=4'h8;
LUT2 \top/processor/n10584_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [232]),
	.F(\top/processor/n10584_15 )
);
defparam \top/processor/n10584_s10 .INIT=4'h8;
LUT2 \top/processor/n10581_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [235]),
	.F(\top/processor/n10581_15 )
);
defparam \top/processor/n10581_s10 .INIT=4'h8;
LUT2 \top/processor/n10580_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [236]),
	.F(\top/processor/n10580_15 )
);
defparam \top/processor/n10580_s10 .INIT=4'h8;
LUT2 \top/processor/n10575_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [241]),
	.F(\top/processor/n10575_15 )
);
defparam \top/processor/n10575_s10 .INIT=4'h8;
LUT2 \top/processor/n10574_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [242]),
	.F(\top/processor/n10574_15 )
);
defparam \top/processor/n10574_s10 .INIT=4'h8;
LUT2 \top/processor/n10572_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [244]),
	.F(\top/processor/n10572_15 )
);
defparam \top/processor/n10572_s10 .INIT=4'h8;
LUT2 \top/processor/n10571_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [245]),
	.F(\top/processor/n10571_15 )
);
defparam \top/processor/n10571_s10 .INIT=4'h8;
LUT2 \top/processor/n10570_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [246]),
	.F(\top/processor/n10570_15 )
);
defparam \top/processor/n10570_s10 .INIT=4'h8;
LUT2 \top/processor/n10569_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [247]),
	.F(\top/processor/n10569_15 )
);
defparam \top/processor/n10569_s10 .INIT=4'h8;
LUT2 \top/processor/n10568_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [248]),
	.F(\top/processor/n10568_15 )
);
defparam \top/processor/n10568_s10 .INIT=4'h8;
LUT2 \top/processor/n10566_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [250]),
	.F(\top/processor/n10566_15 )
);
defparam \top/processor/n10566_s10 .INIT=4'h8;
LUT2 \top/processor/n10564_s10  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [252]),
	.F(\top/processor/n10564_15 )
);
defparam \top/processor/n10564_s10 .INIT=4'h8;
LUT2 \top/processor/n10561_s11  (
	.I0(\top/state_0 [1]),
	.I1(\top/processor/core_hash_out [255]),
	.F(\top/processor/n10561_16 )
);
defparam \top/processor/n10561_s11 .INIT=4'h8;
LUT3 \top/processor/n9789_s11  (
	.I0(\top/state_0 [2]),
	.I1(\top/processor/core_busy ),
	.I2(\top/processor/block_ready ),
	.F(\top/processor/n9789_16 )
);
defparam \top/processor/n9789_s11 .INIT=8'h10;
LUT2 \top/processor/n8408_s2  (
	.I0(\top/processor/core_ready_prev ),
	.I1(\top/processor/core_ready ),
	.F(\top/processor/n8408_6 )
);
defparam \top/processor/n8408_s2 .INIT=4'hB;
LUT2 \top/processor/n10816_s11  (
	.I0(\top/processor/core_hash_out [0]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10816_16 )
);
defparam \top/processor/n10816_s11 .INIT=4'hB;
LUT2 \top/processor/n10813_s11  (
	.I0(\top/processor/core_hash_out [3]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10813_16 )
);
defparam \top/processor/n10813_s11 .INIT=4'hB;
LUT2 \top/processor/n10812_s11  (
	.I0(\top/processor/core_hash_out [4]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10812_16 )
);
defparam \top/processor/n10812_s11 .INIT=4'hB;
LUT2 \top/processor/n10808_s11  (
	.I0(\top/processor/core_hash_out [8]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10808_16 )
);
defparam \top/processor/n10808_s11 .INIT=4'hB;
LUT2 \top/processor/n10806_s11  (
	.I0(\top/processor/core_hash_out [10]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10806_16 )
);
defparam \top/processor/n10806_s11 .INIT=4'hB;
LUT2 \top/processor/n10805_s11  (
	.I0(\top/processor/core_hash_out [11]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10805_16 )
);
defparam \top/processor/n10805_s11 .INIT=4'hB;
LUT2 \top/processor/n10802_s11  (
	.I0(\top/processor/core_hash_out [14]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10802_16 )
);
defparam \top/processor/n10802_s11 .INIT=4'hB;
LUT2 \top/processor/n10801_s11  (
	.I0(\top/processor/core_hash_out [15]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10801_16 )
);
defparam \top/processor/n10801_s11 .INIT=4'hB;
LUT2 \top/processor/n10795_s11  (
	.I0(\top/processor/core_hash_out [21]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10795_16 )
);
defparam \top/processor/n10795_s11 .INIT=4'hB;
LUT2 \top/processor/n10794_s11  (
	.I0(\top/processor/core_hash_out [22]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10794_16 )
);
defparam \top/processor/n10794_s11 .INIT=4'hB;
LUT2 \top/processor/n10793_s11  (
	.I0(\top/processor/core_hash_out [23]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10793_16 )
);
defparam \top/processor/n10793_s11 .INIT=4'hB;
LUT2 \top/processor/n10792_s11  (
	.I0(\top/processor/core_hash_out [24]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10792_16 )
);
defparam \top/processor/n10792_s11 .INIT=4'hB;
LUT2 \top/processor/n10791_s11  (
	.I0(\top/processor/core_hash_out [25]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10791_16 )
);
defparam \top/processor/n10791_s11 .INIT=4'hB;
LUT2 \top/processor/n10789_s11  (
	.I0(\top/processor/core_hash_out [27]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10789_16 )
);
defparam \top/processor/n10789_s11 .INIT=4'hB;
LUT2 \top/processor/n10788_s11  (
	.I0(\top/processor/core_hash_out [28]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10788_16 )
);
defparam \top/processor/n10788_s11 .INIT=4'hB;
LUT2 \top/processor/n10786_s11  (
	.I0(\top/processor/core_hash_out [30]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10786_16 )
);
defparam \top/processor/n10786_s11 .INIT=4'hB;
LUT2 \top/processor/n10784_s11  (
	.I0(\top/processor/core_hash_out [32]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10784_16 )
);
defparam \top/processor/n10784_s11 .INIT=4'hB;
LUT2 \top/processor/n10783_s11  (
	.I0(\top/processor/core_hash_out [33]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10783_16 )
);
defparam \top/processor/n10783_s11 .INIT=4'hB;
LUT2 \top/processor/n10781_s11  (
	.I0(\top/processor/core_hash_out [35]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10781_16 )
);
defparam \top/processor/n10781_s11 .INIT=4'hB;
LUT2 \top/processor/n10779_s11  (
	.I0(\top/processor/core_hash_out [37]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10779_16 )
);
defparam \top/processor/n10779_s11 .INIT=4'hB;
LUT2 \top/processor/n10777_s11  (
	.I0(\top/processor/core_hash_out [39]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10777_16 )
);
defparam \top/processor/n10777_s11 .INIT=4'hB;
LUT2 \top/processor/n10776_s11  (
	.I0(\top/processor/core_hash_out [40]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10776_16 )
);
defparam \top/processor/n10776_s11 .INIT=4'hB;
LUT2 \top/processor/n10773_s11  (
	.I0(\top/processor/core_hash_out [43]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10773_16 )
);
defparam \top/processor/n10773_s11 .INIT=4'hB;
LUT2 \top/processor/n10772_s11  (
	.I0(\top/processor/core_hash_out [44]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10772_16 )
);
defparam \top/processor/n10772_s11 .INIT=4'hB;
LUT2 \top/processor/n10770_s11  (
	.I0(\top/processor/core_hash_out [46]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10770_16 )
);
defparam \top/processor/n10770_s11 .INIT=4'hB;
LUT2 \top/processor/n10769_s11  (
	.I0(\top/processor/core_hash_out [47]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10769_16 )
);
defparam \top/processor/n10769_s11 .INIT=4'hB;
LUT2 \top/processor/n10768_s11  (
	.I0(\top/processor/core_hash_out [48]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10768_16 )
);
defparam \top/processor/n10768_s11 .INIT=4'hB;
LUT2 \top/processor/n10767_s11  (
	.I0(\top/processor/core_hash_out [49]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10767_16 )
);
defparam \top/processor/n10767_s11 .INIT=4'hB;
LUT2 \top/processor/n10761_s11  (
	.I0(\top/processor/core_hash_out [55]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10761_16 )
);
defparam \top/processor/n10761_s11 .INIT=4'hB;
LUT2 \top/processor/n10760_s11  (
	.I0(\top/processor/core_hash_out [56]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10760_16 )
);
defparam \top/processor/n10760_s11 .INIT=4'hB;
LUT2 \top/processor/n10759_s11  (
	.I0(\top/processor/core_hash_out [57]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10759_16 )
);
defparam \top/processor/n10759_s11 .INIT=4'hB;
LUT2 \top/processor/n10758_s11  (
	.I0(\top/processor/core_hash_out [58]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10758_16 )
);
defparam \top/processor/n10758_s11 .INIT=4'hB;
LUT2 \top/processor/n10757_s11  (
	.I0(\top/processor/core_hash_out [59]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10757_16 )
);
defparam \top/processor/n10757_s11 .INIT=4'hB;
LUT2 \top/processor/n10756_s11  (
	.I0(\top/processor/core_hash_out [60]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10756_16 )
);
defparam \top/processor/n10756_s11 .INIT=4'hB;
LUT2 \top/processor/n10750_s11  (
	.I0(\top/processor/core_hash_out [66]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10750_16 )
);
defparam \top/processor/n10750_s11 .INIT=4'hB;
LUT2 \top/processor/n10749_s11  (
	.I0(\top/processor/core_hash_out [67]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10749_16 )
);
defparam \top/processor/n10749_s11 .INIT=4'hB;
LUT2 \top/processor/n10745_s11  (
	.I0(\top/processor/core_hash_out [71]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10745_16 )
);
defparam \top/processor/n10745_s11 .INIT=4'hB;
LUT2 \top/processor/n10741_s11  (
	.I0(\top/processor/core_hash_out [75]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10741_16 )
);
defparam \top/processor/n10741_s11 .INIT=4'hB;
LUT2 \top/processor/n10739_s11  (
	.I0(\top/processor/core_hash_out [77]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10739_16 )
);
defparam \top/processor/n10739_s11 .INIT=4'hB;
LUT2 \top/processor/n10738_s11  (
	.I0(\top/processor/core_hash_out [78]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10738_16 )
);
defparam \top/processor/n10738_s11 .INIT=4'hB;
LUT2 \top/processor/n10736_s11  (
	.I0(\top/processor/core_hash_out [80]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10736_16 )
);
defparam \top/processor/n10736_s11 .INIT=4'hB;
LUT2 \top/processor/n10734_s11  (
	.I0(\top/processor/core_hash_out [82]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10734_16 )
);
defparam \top/processor/n10734_s11 .INIT=4'hB;
LUT2 \top/processor/n10728_s11  (
	.I0(\top/processor/core_hash_out [88]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10728_16 )
);
defparam \top/processor/n10728_s11 .INIT=4'hB;
LUT2 \top/processor/n10727_s11  (
	.I0(\top/processor/core_hash_out [89]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10727_16 )
);
defparam \top/processor/n10727_s11 .INIT=4'hB;
LUT2 \top/processor/n10725_s11  (
	.I0(\top/processor/core_hash_out [91]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10725_16 )
);
defparam \top/processor/n10725_s11 .INIT=4'hB;
LUT2 \top/processor/n10724_s11  (
	.I0(\top/processor/core_hash_out [92]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10724_16 )
);
defparam \top/processor/n10724_s11 .INIT=4'hB;
LUT2 \top/processor/n10721_s11  (
	.I0(\top/processor/core_hash_out [95]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10721_16 )
);
defparam \top/processor/n10721_s11 .INIT=4'hB;
LUT2 \top/processor/n10720_s11  (
	.I0(\top/processor/core_hash_out [96]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10720_16 )
);
defparam \top/processor/n10720_s11 .INIT=4'hB;
LUT2 \top/processor/n10719_s11  (
	.I0(\top/processor/core_hash_out [97]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10719_16 )
);
defparam \top/processor/n10719_s11 .INIT=4'hB;
LUT2 \top/processor/n10718_s11  (
	.I0(\top/processor/core_hash_out [98]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10718_16 )
);
defparam \top/processor/n10718_s11 .INIT=4'hB;
LUT2 \top/processor/n10717_s11  (
	.I0(\top/processor/core_hash_out [99]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10717_16 )
);
defparam \top/processor/n10717_s11 .INIT=4'hB;
LUT2 \top/processor/n10716_s11  (
	.I0(\top/processor/core_hash_out [100]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10716_16 )
);
defparam \top/processor/n10716_s11 .INIT=4'hB;
LUT2 \top/processor/n10715_s11  (
	.I0(\top/processor/core_hash_out [101]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10715_16 )
);
defparam \top/processor/n10715_s11 .INIT=4'hB;
LUT2 \top/processor/n10714_s11  (
	.I0(\top/processor/core_hash_out [102]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10714_16 )
);
defparam \top/processor/n10714_s11 .INIT=4'hB;
LUT2 \top/processor/n10711_s11  (
	.I0(\top/processor/core_hash_out [105]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10711_16 )
);
defparam \top/processor/n10711_s11 .INIT=4'hB;
LUT2 \top/processor/n10708_s11  (
	.I0(\top/processor/core_hash_out [108]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10708_16 )
);
defparam \top/processor/n10708_s11 .INIT=4'hB;
LUT2 \top/processor/n10706_s11  (
	.I0(\top/processor/core_hash_out [110]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10706_16 )
);
defparam \top/processor/n10706_s11 .INIT=4'hB;
LUT2 \top/processor/n10703_s11  (
	.I0(\top/processor/core_hash_out [113]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10703_16 )
);
defparam \top/processor/n10703_s11 .INIT=4'hB;
LUT2 \top/processor/n10702_s11  (
	.I0(\top/processor/core_hash_out [114]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10702_16 )
);
defparam \top/processor/n10702_s11 .INIT=4'hB;
LUT2 \top/processor/n10701_s11  (
	.I0(\top/processor/core_hash_out [115]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10701_16 )
);
defparam \top/processor/n10701_s11 .INIT=4'hB;
LUT2 \top/processor/n10696_s11  (
	.I0(\top/processor/core_hash_out [120]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10696_16 )
);
defparam \top/processor/n10696_s11 .INIT=4'hB;
LUT2 \top/processor/n10692_s11  (
	.I0(\top/processor/core_hash_out [124]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10692_16 )
);
defparam \top/processor/n10692_s11 .INIT=4'hB;
LUT2 \top/processor/n10690_s11  (
	.I0(\top/processor/core_hash_out [126]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10690_16 )
);
defparam \top/processor/n10690_s11 .INIT=4'hB;
LUT2 \top/processor/n10687_s11  (
	.I0(\top/processor/core_hash_out [129]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10687_16 )
);
defparam \top/processor/n10687_s11 .INIT=4'hB;
LUT2 \top/processor/n10685_s11  (
	.I0(\top/processor/core_hash_out [131]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10685_16 )
);
defparam \top/processor/n10685_s11 .INIT=4'hB;
LUT2 \top/processor/n10684_s11  (
	.I0(\top/processor/core_hash_out [132]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10684_16 )
);
defparam \top/processor/n10684_s11 .INIT=4'hB;
LUT2 \top/processor/n10683_s11  (
	.I0(\top/processor/core_hash_out [133]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10683_16 )
);
defparam \top/processor/n10683_s11 .INIT=4'hB;
LUT2 \top/processor/n10680_s11  (
	.I0(\top/processor/core_hash_out [136]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10680_16 )
);
defparam \top/processor/n10680_s11 .INIT=4'hB;
LUT2 \top/processor/n10678_s11  (
	.I0(\top/processor/core_hash_out [138]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10678_16 )
);
defparam \top/processor/n10678_s11 .INIT=4'hB;
LUT2 \top/processor/n10676_s11  (
	.I0(\top/processor/core_hash_out [140]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10676_16 )
);
defparam \top/processor/n10676_s11 .INIT=4'hB;
LUT2 \top/processor/n10675_s11  (
	.I0(\top/processor/core_hash_out [141]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10675_16 )
);
defparam \top/processor/n10675_s11 .INIT=4'hB;
LUT2 \top/processor/n10674_s11  (
	.I0(\top/processor/core_hash_out [142]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10674_16 )
);
defparam \top/processor/n10674_s11 .INIT=4'hB;
LUT2 \top/processor/n10673_s11  (
	.I0(\top/processor/core_hash_out [143]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10673_16 )
);
defparam \top/processor/n10673_s11 .INIT=4'hB;
LUT2 \top/processor/n10672_s11  (
	.I0(\top/processor/core_hash_out [144]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10672_16 )
);
defparam \top/processor/n10672_s11 .INIT=4'hB;
LUT2 \top/processor/n10671_s11  (
	.I0(\top/processor/core_hash_out [145]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10671_16 )
);
defparam \top/processor/n10671_s11 .INIT=4'hB;
LUT2 \top/processor/n10670_s11  (
	.I0(\top/processor/core_hash_out [146]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10670_16 )
);
defparam \top/processor/n10670_s11 .INIT=4'hB;
LUT2 \top/processor/n10669_s11  (
	.I0(\top/processor/core_hash_out [147]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10669_16 )
);
defparam \top/processor/n10669_s11 .INIT=4'hB;
LUT2 \top/processor/n10666_s11  (
	.I0(\top/processor/core_hash_out [150]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10666_16 )
);
defparam \top/processor/n10666_s11 .INIT=4'hB;
LUT2 \top/processor/n10664_s11  (
	.I0(\top/processor/core_hash_out [152]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10664_16 )
);
defparam \top/processor/n10664_s11 .INIT=4'hB;
LUT2 \top/processor/n10662_s11  (
	.I0(\top/processor/core_hash_out [154]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10662_16 )
);
defparam \top/processor/n10662_s11 .INIT=4'hB;
LUT2 \top/processor/n10659_s11  (
	.I0(\top/processor/core_hash_out [157]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10659_16 )
);
defparam \top/processor/n10659_s11 .INIT=4'hB;
LUT2 \top/processor/n10657_s11  (
	.I0(\top/processor/core_hash_out [159]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10657_16 )
);
defparam \top/processor/n10657_s11 .INIT=4'hB;
LUT2 \top/processor/n10655_s11  (
	.I0(\top/processor/core_hash_out [161]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10655_16 )
);
defparam \top/processor/n10655_s11 .INIT=4'hB;
LUT2 \top/processor/n10652_s11  (
	.I0(\top/processor/core_hash_out [164]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10652_16 )
);
defparam \top/processor/n10652_s11 .INIT=4'hB;
LUT2 \top/processor/n10651_s11  (
	.I0(\top/processor/core_hash_out [165]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10651_16 )
);
defparam \top/processor/n10651_s11 .INIT=4'hB;
LUT2 \top/processor/n10650_s11  (
	.I0(\top/processor/core_hash_out [166]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10650_16 )
);
defparam \top/processor/n10650_s11 .INIT=4'hB;
LUT2 \top/processor/n10648_s11  (
	.I0(\top/processor/core_hash_out [168]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10648_16 )
);
defparam \top/processor/n10648_s11 .INIT=4'hB;
LUT2 \top/processor/n10647_s11  (
	.I0(\top/processor/core_hash_out [169]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10647_16 )
);
defparam \top/processor/n10647_s11 .INIT=4'hB;
LUT2 \top/processor/n10644_s11  (
	.I0(\top/processor/core_hash_out [172]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10644_16 )
);
defparam \top/processor/n10644_s11 .INIT=4'hB;
LUT2 \top/processor/n10643_s11  (
	.I0(\top/processor/core_hash_out [173]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10643_16 )
);
defparam \top/processor/n10643_s11 .INIT=4'hB;
LUT2 \top/processor/n10642_s11  (
	.I0(\top/processor/core_hash_out [174]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10642_16 )
);
defparam \top/processor/n10642_s11 .INIT=4'hB;
LUT2 \top/processor/n10641_s11  (
	.I0(\top/processor/core_hash_out [175]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10641_16 )
);
defparam \top/processor/n10641_s11 .INIT=4'hB;
LUT2 \top/processor/n10639_s11  (
	.I0(\top/processor/core_hash_out [177]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10639_16 )
);
defparam \top/processor/n10639_s11 .INIT=4'hB;
LUT2 \top/processor/n10638_s11  (
	.I0(\top/processor/core_hash_out [178]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10638_16 )
);
defparam \top/processor/n10638_s11 .INIT=4'hB;
LUT2 \top/processor/n10637_s11  (
	.I0(\top/processor/core_hash_out [179]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10637_16 )
);
defparam \top/processor/n10637_s11 .INIT=4'hB;
LUT2 \top/processor/n10635_s11  (
	.I0(\top/processor/core_hash_out [181]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10635_16 )
);
defparam \top/processor/n10635_s11 .INIT=4'hB;
LUT2 \top/processor/n10634_s11  (
	.I0(\top/processor/core_hash_out [182]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10634_16 )
);
defparam \top/processor/n10634_s11 .INIT=4'hB;
LUT2 \top/processor/n10630_s11  (
	.I0(\top/processor/core_hash_out [186]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10630_16 )
);
defparam \top/processor/n10630_s11 .INIT=4'hB;
LUT2 \top/processor/n10629_s11  (
	.I0(\top/processor/core_hash_out [187]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10629_16 )
);
defparam \top/processor/n10629_s11 .INIT=4'hB;
LUT2 \top/processor/n10628_s11  (
	.I0(\top/processor/core_hash_out [188]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10628_16 )
);
defparam \top/processor/n10628_s11 .INIT=4'hB;
LUT2 \top/processor/n10627_s11  (
	.I0(\top/processor/core_hash_out [189]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10627_16 )
);
defparam \top/processor/n10627_s11 .INIT=4'hB;
LUT2 \top/processor/n10624_s11  (
	.I0(\top/processor/core_hash_out [192]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10624_16 )
);
defparam \top/processor/n10624_s11 .INIT=4'hB;
LUT2 \top/processor/n10622_s11  (
	.I0(\top/processor/core_hash_out [194]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10622_16 )
);
defparam \top/processor/n10622_s11 .INIT=4'hB;
LUT2 \top/processor/n10617_s11  (
	.I0(\top/processor/core_hash_out [199]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10617_16 )
);
defparam \top/processor/n10617_s11 .INIT=4'hB;
LUT2 \top/processor/n10615_s11  (
	.I0(\top/processor/core_hash_out [201]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10615_16 )
);
defparam \top/processor/n10615_s11 .INIT=4'hB;
LUT2 \top/processor/n10614_s11  (
	.I0(\top/processor/core_hash_out [202]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10614_16 )
);
defparam \top/processor/n10614_s11 .INIT=4'hB;
LUT2 \top/processor/n10613_s11  (
	.I0(\top/processor/core_hash_out [203]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10613_16 )
);
defparam \top/processor/n10613_s11 .INIT=4'hB;
LUT2 \top/processor/n10611_s11  (
	.I0(\top/processor/core_hash_out [205]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10611_16 )
);
defparam \top/processor/n10611_s11 .INIT=4'hB;
LUT2 \top/processor/n10609_s11  (
	.I0(\top/processor/core_hash_out [207]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10609_16 )
);
defparam \top/processor/n10609_s11 .INIT=4'hB;
LUT2 \top/processor/n10608_s11  (
	.I0(\top/processor/core_hash_out [208]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10608_16 )
);
defparam \top/processor/n10608_s11 .INIT=4'hB;
LUT2 \top/processor/n10607_s11  (
	.I0(\top/processor/core_hash_out [209]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10607_16 )
);
defparam \top/processor/n10607_s11 .INIT=4'hB;
LUT2 \top/processor/n10606_s11  (
	.I0(\top/processor/core_hash_out [210]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10606_16 )
);
defparam \top/processor/n10606_s11 .INIT=4'hB;
LUT2 \top/processor/n10603_s11  (
	.I0(\top/processor/core_hash_out [213]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10603_16 )
);
defparam \top/processor/n10603_s11 .INIT=4'hB;
LUT2 \top/processor/n10602_s11  (
	.I0(\top/processor/core_hash_out [214]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10602_16 )
);
defparam \top/processor/n10602_s11 .INIT=4'hB;
LUT2 \top/processor/n10600_s11  (
	.I0(\top/processor/core_hash_out [216]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10600_16 )
);
defparam \top/processor/n10600_s11 .INIT=4'hB;
LUT2 \top/processor/n10599_s11  (
	.I0(\top/processor/core_hash_out [217]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10599_16 )
);
defparam \top/processor/n10599_s11 .INIT=4'hB;
LUT2 \top/processor/n10597_s11  (
	.I0(\top/processor/core_hash_out [219]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10597_16 )
);
defparam \top/processor/n10597_s11 .INIT=4'hB;
LUT2 \top/processor/n10596_s11  (
	.I0(\top/processor/core_hash_out [220]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10596_16 )
);
defparam \top/processor/n10596_s11 .INIT=4'hB;
LUT2 \top/processor/n10595_s11  (
	.I0(\top/processor/core_hash_out [221]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10595_16 )
);
defparam \top/processor/n10595_s11 .INIT=4'hB;
LUT2 \top/processor/n10593_s11  (
	.I0(\top/processor/core_hash_out [223]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10593_16 )
);
defparam \top/processor/n10593_s11 .INIT=4'hB;
LUT2 \top/processor/n10592_s11  (
	.I0(\top/processor/core_hash_out [224]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10592_16 )
);
defparam \top/processor/n10592_s11 .INIT=4'hB;
LUT2 \top/processor/n10591_s11  (
	.I0(\top/processor/core_hash_out [225]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10591_16 )
);
defparam \top/processor/n10591_s11 .INIT=4'hB;
LUT2 \top/processor/n10590_s11  (
	.I0(\top/processor/core_hash_out [226]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10590_16 )
);
defparam \top/processor/n10590_s11 .INIT=4'hB;
LUT2 \top/processor/n10587_s11  (
	.I0(\top/processor/core_hash_out [229]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10587_16 )
);
defparam \top/processor/n10587_s11 .INIT=4'hB;
LUT2 \top/processor/n10586_s11  (
	.I0(\top/processor/core_hash_out [230]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10586_16 )
);
defparam \top/processor/n10586_s11 .INIT=4'hB;
LUT2 \top/processor/n10583_s11  (
	.I0(\top/processor/core_hash_out [233]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10583_16 )
);
defparam \top/processor/n10583_s11 .INIT=4'hB;
LUT2 \top/processor/n10582_s11  (
	.I0(\top/processor/core_hash_out [234]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10582_16 )
);
defparam \top/processor/n10582_s11 .INIT=4'hB;
LUT2 \top/processor/n10579_s11  (
	.I0(\top/processor/core_hash_out [237]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10579_16 )
);
defparam \top/processor/n10579_s11 .INIT=4'hB;
LUT2 \top/processor/n10578_s11  (
	.I0(\top/processor/core_hash_out [238]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10578_16 )
);
defparam \top/processor/n10578_s11 .INIT=4'hB;
LUT2 \top/processor/n10577_s11  (
	.I0(\top/processor/core_hash_out [239]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10577_16 )
);
defparam \top/processor/n10577_s11 .INIT=4'hB;
LUT2 \top/processor/n10576_s11  (
	.I0(\top/processor/core_hash_out [240]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10576_16 )
);
defparam \top/processor/n10576_s11 .INIT=4'hB;
LUT2 \top/processor/n10573_s11  (
	.I0(\top/processor/core_hash_out [243]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10573_16 )
);
defparam \top/processor/n10573_s11 .INIT=4'hB;
LUT2 \top/processor/n10567_s11  (
	.I0(\top/processor/core_hash_out [249]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10567_16 )
);
defparam \top/processor/n10567_s11 .INIT=4'hB;
LUT2 \top/processor/n10565_s11  (
	.I0(\top/processor/core_hash_out [251]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10565_16 )
);
defparam \top/processor/n10565_s11 .INIT=4'hB;
LUT2 \top/processor/n10563_s11  (
	.I0(\top/processor/core_hash_out [253]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10563_16 )
);
defparam \top/processor/n10563_s11 .INIT=4'hB;
LUT2 \top/processor/n10562_s11  (
	.I0(\top/processor/core_hash_out [254]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n10562_16 )
);
defparam \top/processor/n10562_s11 .INIT=4'hB;
LUT2 \top/processor/n9790_s6  (
	.I0(\top/state_0 [0]),
	.I1(\top/state_0 [1]),
	.F(\top/processor/n9790_11 )
);
defparam \top/processor/n9790_s6 .INIT=4'h8;
LUT4 \top/processor/n10817_s10  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [4]),
	.I2(\top/processor/pad_index [5]),
	.I3(\top/processor/block_buffer_63_10 ),
	.F(\top/processor/n10817_15 )
);
defparam \top/processor/n10817_s10 .INIT=16'h0100;
LUT2 \top/processor/n11265_s9  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/n11374_20 ),
	.F(\top/processor/n11265_13 )
);
defparam \top/processor/n11265_s9 .INIT=4'h1;
LUT3 \top/processor/n11361_s11  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [3]),
	.I2(\top/processor/byte_index [5]),
	.F(\top/processor/n11361_17 )
);
defparam \top/processor/n11361_s11 .INIT=8'h80;
LUT4 \top/processor/n11364_s22  (
	.I0(\top/processor/n7631_12 ),
	.I1(\top/data_last ),
	.I2(\top/data_valid ),
	.I3(\top/processor/n11370_19 ),
	.F(\top/processor/n11364_28 )
);
defparam \top/processor/n11364_s22 .INIT=16'h4F00;
LUT4 \top/processor/n11362_s11  (
	.I0(\top/processor/n8408_6 ),
	.I1(\top/processor/n11362_19 ),
	.I2(\top/processor/n11374_20 ),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11362_18 )
);
defparam \top/processor/n11362_s11 .INIT=16'hEE0F;
LUT4 \top/processor/state_1_s5  (
	.I0(\top/processor/n7631_12 ),
	.I1(\top/processor/state_1_10 ),
	.I2(\top/state_0 [0]),
	.I3(\top/data_valid ),
	.F(\top/processor/state_1_9 )
);
defparam \top/processor/state_1_s5 .INIT=16'hE33C;
LUT3 \top/processor/hash_state_255_s5  (
	.I0(\top/state_0 [0]),
	.I1(\top/state_0 [1]),
	.I2(\top/data_last ),
	.F(\top/processor/hash_state_255_8 )
);
defparam \top/processor/hash_state_255_s5 .INIT=8'h10;
LUT2 \top/processor/seen_last_s5  (
	.I0(\top/data_valid ),
	.I1(\top/state_0 [0]),
	.F(\top/processor/seen_last_9 )
);
defparam \top/processor/seen_last_s5 .INIT=4'h4;
LUT4 \top/processor/need_length_block_s5  (
	.I0(\top/data_valid ),
	.I1(\top/processor/n7631_12 ),
	.I2(\top/state_0 [0]),
	.I3(\top/data_last ),
	.F(\top/processor/need_length_block_9 )
);
defparam \top/processor/need_length_block_s5 .INIT=16'h8F00;
LUT4 \top/processor/need_length_block_s6  (
	.I0(\top/state_0 [0]),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/n10817_15 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/need_length_block_10 )
);
defparam \top/processor/need_length_block_s6 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_511_s5  (
	.I0(\top/processor/n8408_6 ),
	.I1(\top/processor/need_length_block ),
	.I2(\top/processor/seen_last ),
	.I3(\top/processor/n9790_11 ),
	.F(\top/processor/block_buffer_511_9 )
);
defparam \top/processor/block_buffer_511_s5 .INIT=16'h4000;
LUT3 \top/processor/block_buffer_511_s6  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_319_9 ),
	.I2(\top/processor/block_buffer_511_13 ),
	.F(\top/processor/block_buffer_511_10 )
);
defparam \top/processor/block_buffer_511_s6 .INIT=8'h40;
LUT2 \top/processor/block_buffer_511_s7  (
	.I0(\top/state_0 [2]),
	.I1(rst),
	.F(\top/processor/block_buffer_511_11 )
);
defparam \top/processor/block_buffer_511_s7 .INIT=4'h1;
LUT4 \top/processor/block_buffer_503_s5  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [4]),
	.I2(\top/processor/pad_index [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/block_buffer_503_9 )
);
defparam \top/processor/block_buffer_503_s5 .INIT=16'h0100;
LUT4 \top/processor/block_buffer_503_s6  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [2]),
	.I3(\top/processor/pad_index [0]),
	.F(\top/processor/block_buffer_503_10 )
);
defparam \top/processor/block_buffer_503_s6 .INIT=16'h0100;
LUT4 \top/processor/block_buffer_503_s7  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_511_13 ),
	.I2(\top/processor/block_buffer_439_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_503_11 )
);
defparam \top/processor/block_buffer_503_s7 .INIT=16'h00BF;
LUT3 \top/processor/block_buffer_495_s5  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/pad_index [2]),
	.I2(\top/processor/pad_index [1]),
	.F(\top/processor/block_buffer_495_9 )
);
defparam \top/processor/block_buffer_495_s5 .INIT=8'h10;
LUT4 \top/processor/block_buffer_495_s7  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_511_13 ),
	.I2(\top/processor/block_buffer_431_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_495_11 )
);
defparam \top/processor/block_buffer_495_s7 .INIT=16'h00BF;
LUT3 \top/processor/block_buffer_487_s5  (
	.I0(\top/processor/pad_index [2]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [0]),
	.F(\top/processor/block_buffer_487_9 )
);
defparam \top/processor/block_buffer_487_s5 .INIT=8'h40;
LUT4 \top/processor/block_buffer_487_s6  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_511_13 ),
	.I2(\top/processor/block_buffer_423_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_487_10 )
);
defparam \top/processor/block_buffer_487_s6 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_479_s5  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [1]),
	.I3(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_479_9 )
);
defparam \top/processor/block_buffer_479_s5 .INIT=16'h0100;
LUT4 \top/processor/block_buffer_479_s6  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_511_13 ),
	.I2(\top/processor/block_buffer_415_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_479_10 )
);
defparam \top/processor/block_buffer_479_s6 .INIT=16'h00BF;
LUT3 \top/processor/block_buffer_471_s5  (
	.I0(\top/processor/pad_index [1]),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_471_9 )
);
defparam \top/processor/block_buffer_471_s5 .INIT=8'h40;
LUT4 \top/processor/block_buffer_471_s6  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_511_13 ),
	.I2(\top/processor/block_buffer_407_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_471_10 )
);
defparam \top/processor/block_buffer_471_s6 .INIT=16'h00BF;
LUT3 \top/processor/block_buffer_463_s5  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_463_9 )
);
defparam \top/processor/block_buffer_463_s5 .INIT=8'h40;
LUT4 \top/processor/block_buffer_463_s6  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_511_13 ),
	.I2(\top/processor/block_buffer_399_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_463_10 )
);
defparam \top/processor/block_buffer_463_s6 .INIT=16'h00BF;
LUT3 \top/processor/block_buffer_455_s5  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_455_9 )
);
defparam \top/processor/block_buffer_455_s5 .INIT=8'h80;
LUT4 \top/processor/block_buffer_455_s6  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/block_buffer_391_9 ),
	.I2(\top/processor/block_buffer_511_13 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_455_10 )
);
defparam \top/processor/block_buffer_455_s6 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_447_s5  (
	.I0(\top/processor/n7631_8 ),
	.I1(\top/processor/block_buffer_447_10 ),
	.I2(\top/processor/block_buffer_447_11 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_447_9 )
);
defparam \top/processor/block_buffer_447_s5 .INIT=16'h0007;
LUT3 \top/processor/block_buffer_439_s5  (
	.I0(\top/processor/byte_index [1]),
	.I1(\top/processor/byte_index [2]),
	.I2(\top/processor/byte_index [0]),
	.F(\top/processor/block_buffer_439_9 )
);
defparam \top/processor/block_buffer_439_s5 .INIT=8'h10;
LUT4 \top/processor/block_buffer_439_s6  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [5]),
	.I2(\top/processor/block_buffer_511_12 ),
	.I3(\top/processor/byte_index [3]),
	.F(\top/processor/block_buffer_439_10 )
);
defparam \top/processor/block_buffer_439_s6 .INIT=16'h0100;
LUT3 \top/processor/block_buffer_439_s7  (
	.I0(\top/processor/block_buffer_439_12 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_439_11 )
);
defparam \top/processor/block_buffer_439_s7 .INIT=8'h07;
LUT3 \top/processor/block_buffer_431_s5  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [2]),
	.I2(\top/processor/byte_index [1]),
	.F(\top/processor/block_buffer_431_9 )
);
defparam \top/processor/block_buffer_431_s5 .INIT=8'h10;
LUT3 \top/processor/block_buffer_431_s6  (
	.I0(\top/processor/block_buffer_431_13 ),
	.I1(\top/processor/block_buffer_439_12 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_431_10 )
);
defparam \top/processor/block_buffer_431_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_423_s5  (
	.I0(\top/processor/byte_index [2]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [0]),
	.F(\top/processor/block_buffer_423_9 )
);
defparam \top/processor/block_buffer_423_s5 .INIT=8'h40;
LUT3 \top/processor/block_buffer_423_s6  (
	.I0(\top/processor/block_buffer_423_11 ),
	.I1(\top/processor/block_buffer_439_12 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_423_10 )
);
defparam \top/processor/block_buffer_423_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_415_s5  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [2]),
	.F(\top/processor/block_buffer_415_9 )
);
defparam \top/processor/block_buffer_415_s5 .INIT=8'h10;
LUT3 \top/processor/block_buffer_415_s6  (
	.I0(\top/processor/block_buffer_439_12 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_415_10 )
);
defparam \top/processor/block_buffer_415_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_407_s5  (
	.I0(\top/processor/byte_index [1]),
	.I1(\top/processor/byte_index [0]),
	.I2(\top/processor/byte_index [2]),
	.F(\top/processor/block_buffer_407_9 )
);
defparam \top/processor/block_buffer_407_s5 .INIT=8'h40;
LUT3 \top/processor/block_buffer_407_s6  (
	.I0(\top/processor/block_buffer_407_11 ),
	.I1(\top/processor/block_buffer_439_12 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_407_10 )
);
defparam \top/processor/block_buffer_407_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_399_s5  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [2]),
	.F(\top/processor/block_buffer_399_9 )
);
defparam \top/processor/block_buffer_399_s5 .INIT=8'h40;
LUT3 \top/processor/block_buffer_399_s6  (
	.I0(\top/processor/block_buffer_399_13 ),
	.I1(\top/processor/block_buffer_439_12 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_399_10 )
);
defparam \top/processor/block_buffer_399_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_391_s5  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [2]),
	.F(\top/processor/block_buffer_391_9 )
);
defparam \top/processor/block_buffer_391_s5 .INIT=8'h80;
LUT4 \top/processor/block_buffer_391_s6  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_439_12 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_391_10 )
);
defparam \top/processor/block_buffer_391_s6 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_383_s5  (
	.I0(\top/processor/n7631_8 ),
	.I1(\top/processor/pad_index [4]),
	.I2(\top/processor/block_buffer_383_10 ),
	.I3(\top/processor/block_buffer_383_11 ),
	.F(\top/processor/block_buffer_383_9 )
);
defparam \top/processor/block_buffer_383_s5 .INIT=16'hFCA0;
LUT4 \top/processor/block_buffer_375_s5  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/byte_index [5]),
	.I2(\top/processor/block_buffer_511_12 ),
	.I3(\top/processor/byte_index [4]),
	.F(\top/processor/block_buffer_375_9 )
);
defparam \top/processor/block_buffer_375_s5 .INIT=16'h0100;
LUT3 \top/processor/block_buffer_375_s6  (
	.I0(\top/processor/block_buffer_375_11 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_375_10 )
);
defparam \top/processor/block_buffer_375_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_367_s5  (
	.I0(\top/processor/block_buffer_375_11 ),
	.I1(\top/processor/block_buffer_431_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_367_9 )
);
defparam \top/processor/block_buffer_367_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_359_s5  (
	.I0(\top/processor/block_buffer_375_11 ),
	.I1(\top/processor/block_buffer_423_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_359_9 )
);
defparam \top/processor/block_buffer_359_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_351_s5  (
	.I0(\top/processor/block_buffer_375_11 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_351_9 )
);
defparam \top/processor/block_buffer_351_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_343_s5  (
	.I0(\top/processor/block_buffer_375_11 ),
	.I1(\top/processor/block_buffer_407_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_343_9 )
);
defparam \top/processor/block_buffer_343_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_335_s5  (
	.I0(\top/processor/block_buffer_375_11 ),
	.I1(\top/processor/block_buffer_399_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_335_9 )
);
defparam \top/processor/block_buffer_335_s5 .INIT=8'h07;
LUT4 \top/processor/block_buffer_327_s5  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_375_11 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_327_9 )
);
defparam \top/processor/block_buffer_327_s5 .INIT=16'h00BF;
LUT3 \top/processor/block_buffer_319_s5  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [2]),
	.F(\top/processor/block_buffer_319_9 )
);
defparam \top/processor/block_buffer_319_s5 .INIT=8'h01;
LUT4 \top/processor/block_buffer_319_s6  (
	.I0(\top/processor/byte_index [5]),
	.I1(\top/processor/block_buffer_511_12 ),
	.I2(\top/processor/byte_index [4]),
	.I3(\top/processor/byte_index [3]),
	.F(\top/processor/block_buffer_319_10 )
);
defparam \top/processor/block_buffer_319_s6 .INIT=16'h1000;
LUT3 \top/processor/block_buffer_319_s7  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_319_15 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_319_11 )
);
defparam \top/processor/block_buffer_319_s7 .INIT=8'h07;
LUT3 \top/processor/block_buffer_311_s5  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_311_9 )
);
defparam \top/processor/block_buffer_311_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_303_s5  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_431_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_303_9 )
);
defparam \top/processor/block_buffer_303_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_295_s5  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_423_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_295_9 )
);
defparam \top/processor/block_buffer_295_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_287_s5  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_287_9 )
);
defparam \top/processor/block_buffer_287_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_279_s5  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_407_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_279_9 )
);
defparam \top/processor/block_buffer_279_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_271_s5  (
	.I0(\top/processor/block_buffer_319_17 ),
	.I1(\top/processor/block_buffer_399_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_271_9 )
);
defparam \top/processor/block_buffer_271_s5 .INIT=8'h07;
LUT4 \top/processor/block_buffer_263_s5  (
	.I0(\top/processor/pad_index [5]),
	.I1(\top/processor/block_buffer_263_12 ),
	.I2(\top/processor/block_buffer_455_9 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_263_9 )
);
defparam \top/processor/block_buffer_263_s5 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_255_s5  (
	.I0(\top/processor/n7631_8 ),
	.I1(\top/processor/pad_index [5]),
	.I2(\top/processor/block_buffer_255_10 ),
	.I3(\top/processor/block_buffer_255_11 ),
	.F(\top/processor/block_buffer_255_9 )
);
defparam \top/processor/block_buffer_255_s5 .INIT=16'hFCA0;
LUT4 \top/processor/block_buffer_247_s5  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [3]),
	.I2(\top/processor/block_buffer_511_12 ),
	.I3(\top/processor/byte_index [5]),
	.F(\top/processor/block_buffer_247_9 )
);
defparam \top/processor/block_buffer_247_s5 .INIT=16'h0100;
LUT3 \top/processor/block_buffer_247_s6  (
	.I0(\top/processor/block_buffer_247_11 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_247_10 )
);
defparam \top/processor/block_buffer_247_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_239_s5  (
	.I0(\top/processor/block_buffer_247_11 ),
	.I1(\top/processor/block_buffer_431_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_239_9 )
);
defparam \top/processor/block_buffer_239_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_231_s5  (
	.I0(\top/processor/block_buffer_247_11 ),
	.I1(\top/processor/block_buffer_423_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_231_9 )
);
defparam \top/processor/block_buffer_231_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_223_s5  (
	.I0(\top/processor/block_buffer_247_11 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_223_9 )
);
defparam \top/processor/block_buffer_223_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_215_s5  (
	.I0(\top/processor/block_buffer_247_11 ),
	.I1(\top/processor/block_buffer_407_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_215_9 )
);
defparam \top/processor/block_buffer_215_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_207_s5  (
	.I0(\top/processor/block_buffer_247_11 ),
	.I1(\top/processor/block_buffer_399_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_207_9 )
);
defparam \top/processor/block_buffer_207_s5 .INIT=8'h07;
LUT4 \top/processor/block_buffer_199_s5  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_247_11 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_199_9 )
);
defparam \top/processor/block_buffer_199_s5 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_191_s5  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/block_buffer_511_12 ),
	.I2(\top/processor/byte_index [5]),
	.I3(\top/processor/byte_index [3]),
	.F(\top/processor/block_buffer_191_9 )
);
defparam \top/processor/block_buffer_191_s5 .INIT=16'h1000;
LUT3 \top/processor/block_buffer_191_s6  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_319_15 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_191_10 )
);
defparam \top/processor/block_buffer_191_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_183_s5  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_183_9 )
);
defparam \top/processor/block_buffer_183_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_175_s5  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_431_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_175_9 )
);
defparam \top/processor/block_buffer_175_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_167_s5  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_423_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_167_9 )
);
defparam \top/processor/block_buffer_167_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_159_s5  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_159_9 )
);
defparam \top/processor/block_buffer_159_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_151_s5  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_407_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_151_9 )
);
defparam \top/processor/block_buffer_151_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_143_s5  (
	.I0(\top/processor/block_buffer_191_11 ),
	.I1(\top/processor/block_buffer_399_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_143_9 )
);
defparam \top/processor/block_buffer_143_s5 .INIT=8'h07;
LUT4 \top/processor/block_buffer_135_s5  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_191_11 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_135_9 )
);
defparam \top/processor/block_buffer_135_s5 .INIT=16'h00BF;
LUT4 \top/processor/block_buffer_127_s5  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/block_buffer_511_12 ),
	.I2(\top/processor/byte_index [5]),
	.I3(\top/processor/byte_index [4]),
	.F(\top/processor/block_buffer_127_9 )
);
defparam \top/processor/block_buffer_127_s5 .INIT=16'h1000;
LUT3 \top/processor/block_buffer_127_s6  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_319_15 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_127_10 )
);
defparam \top/processor/block_buffer_127_s6 .INIT=8'h07;
LUT3 \top/processor/block_buffer_119_s5  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_503_10 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_119_9 )
);
defparam \top/processor/block_buffer_119_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_111_s5  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_431_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_111_9 )
);
defparam \top/processor/block_buffer_111_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_103_s5  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_423_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_103_9 )
);
defparam \top/processor/block_buffer_103_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_95_s5  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_479_9 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_95_9 )
);
defparam \top/processor/block_buffer_95_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_87_s5  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_407_11 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_87_9 )
);
defparam \top/processor/block_buffer_87_s5 .INIT=8'h07;
LUT3 \top/processor/block_buffer_79_s5  (
	.I0(\top/processor/block_buffer_127_11 ),
	.I1(\top/processor/block_buffer_399_13 ),
	.I2(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_79_9 )
);
defparam \top/processor/block_buffer_79_s5 .INIT=8'h07;
LUT4 \top/processor/block_buffer_71_s5  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_127_11 ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/block_buffer_71_9 )
);
defparam \top/processor/block_buffer_71_s5 .INIT=16'h00BF;
LUT2 \top/processor/block_buffer_63_s5  (
	.I0(\top/processor/pad_index [5]),
	.I1(\top/processor/block_buffer_263_12 ),
	.F(\top/processor/block_buffer_63_9 )
);
defparam \top/processor/block_buffer_63_s5 .INIT=4'h8;
LUT3 \top/processor/block_buffer_63_s6  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_63_10 )
);
defparam \top/processor/block_buffer_63_s6 .INIT=8'h01;
LUT4 \top/processor/block_buffer_63_s7  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_319_9 ),
	.I3(\top/processor/n7631_10 ),
	.F(\top/processor/block_buffer_63_11 )
);
defparam \top/processor/block_buffer_63_s7 .INIT=16'hBF00;
LUT3 \top/processor/block_buffer_55_s5  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_439_9 ),
	.F(\top/processor/block_buffer_55_9 )
);
defparam \top/processor/block_buffer_55_s5 .INIT=8'h40;
LUT4 \top/processor/block_buffer_55_s6  (
	.I0(\top/processor/pad_index [1]),
	.I1(\top/processor/pad_index [2]),
	.I2(\top/processor/pad_index [0]),
	.I3(\top/processor/block_buffer_63_9 ),
	.F(\top/processor/block_buffer_55_10 )
);
defparam \top/processor/block_buffer_55_s6 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_47_s5  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_431_9 ),
	.I3(\top/processor/n7631_10 ),
	.F(\top/processor/block_buffer_47_9 )
);
defparam \top/processor/block_buffer_47_s5 .INIT=16'hBF00;
LUT4 \top/processor/block_buffer_39_s5  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_423_9 ),
	.I3(\top/processor/n7631_10 ),
	.F(\top/processor/block_buffer_39_9 )
);
defparam \top/processor/block_buffer_39_s5 .INIT=16'hBF00;
LUT3 \top/processor/block_buffer_31_s5  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_415_9 ),
	.F(\top/processor/block_buffer_31_9 )
);
defparam \top/processor/block_buffer_31_s5 .INIT=8'h40;
LUT4 \top/processor/block_buffer_31_s6  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [2]),
	.I3(\top/processor/block_buffer_63_9 ),
	.F(\top/processor/block_buffer_31_10 )
);
defparam \top/processor/block_buffer_31_s6 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_23_s5  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_407_9 ),
	.I3(\top/processor/n7631_10 ),
	.F(\top/processor/block_buffer_23_9 )
);
defparam \top/processor/block_buffer_23_s5 .INIT=16'hBF00;
LUT4 \top/processor/block_buffer_15_s5  (
	.I0(\top/processor/block_buffer_511_12 ),
	.I1(\top/processor/n11361_17 ),
	.I2(\top/processor/block_buffer_399_9 ),
	.I3(\top/processor/n7631_10 ),
	.F(\top/processor/block_buffer_15_9 )
);
defparam \top/processor/block_buffer_15_s5 .INIT=16'hBF00;
LUT4 \top/processor/block_buffer_7_s5  (
	.I0(\top/processor/block_buffer_63_9 ),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/block_buffer_511_12 ),
	.I3(\top/processor/n7631_12 ),
	.F(\top/processor/block_buffer_7_9 )
);
defparam \top/processor/block_buffer_7_s5 .INIT=16'h7077;
LUT3 \top/processor/n11435_s10  (
	.I0(\top/processor/total_bits [5]),
	.I1(\top/processor/total_bits [4]),
	.I2(\top/processor/total_bits [3]),
	.F(\top/processor/n11435_15 )
);
defparam \top/processor/n11435_s10 .INIT=8'h80;
LUT4 \top/processor/n11434_s10  (
	.I0(\top/processor/total_bits [6]),
	.I1(\top/processor/total_bits [5]),
	.I2(\top/processor/total_bits [4]),
	.I3(\top/processor/total_bits [3]),
	.F(\top/processor/n11434_15 )
);
defparam \top/processor/n11434_s10 .INIT=16'h8000;
LUT3 \top/processor/n11432_s10  (
	.I0(\top/processor/total_bits [8]),
	.I1(\top/processor/total_bits [7]),
	.I2(\top/processor/n11434_15 ),
	.F(\top/processor/n11432_15 )
);
defparam \top/processor/n11432_s10 .INIT=8'h80;
LUT4 \top/processor/n11431_s10  (
	.I0(\top/processor/total_bits [9]),
	.I1(\top/processor/total_bits [8]),
	.I2(\top/processor/total_bits [7]),
	.I3(\top/processor/n11434_15 ),
	.F(\top/processor/n11431_15 )
);
defparam \top/processor/n11431_s10 .INIT=16'h8000;
LUT2 \top/processor/n11430_s10  (
	.I0(\top/processor/total_bits [10]),
	.I1(\top/processor/n11431_15 ),
	.F(\top/processor/n11430_15 )
);
defparam \top/processor/n11430_s10 .INIT=4'h8;
LUT2 \top/processor/n11428_s10  (
	.I0(\top/processor/total_bits [12]),
	.I1(\top/processor/total_bits [11]),
	.F(\top/processor/n11428_15 )
);
defparam \top/processor/n11428_s10 .INIT=4'h8;
LUT4 \top/processor/n11425_s10  (
	.I0(\top/processor/total_bits [15]),
	.I1(\top/processor/total_bits [14]),
	.I2(\top/processor/total_bits [13]),
	.I3(\top/processor/n11428_15 ),
	.F(\top/processor/n11425_15 )
);
defparam \top/processor/n11425_s10 .INIT=16'h8000;
LUT2 \top/processor/n11423_s10  (
	.I0(\top/processor/total_bits [17]),
	.I1(\top/processor/n11424_17 ),
	.F(\top/processor/n11423_15 )
);
defparam \top/processor/n11423_s10 .INIT=4'h8;
LUT4 \top/processor/n11420_s10  (
	.I0(\top/processor/n11420_16 ),
	.I1(\top/processor/total_bits [20]),
	.I2(\top/processor/total_bits [19]),
	.I3(\top/processor/n11430_15 ),
	.F(\top/processor/n11420_15 )
);
defparam \top/processor/n11420_s10 .INIT=16'h8000;
LUT3 \top/processor/n11418_s10  (
	.I0(\top/processor/total_bits [22]),
	.I1(\top/processor/total_bits [21]),
	.I2(\top/processor/n11420_15 ),
	.F(\top/processor/n11418_15 )
);
defparam \top/processor/n11418_s10 .INIT=8'h80;
LUT3 \top/processor/n11417_s10  (
	.I0(\top/processor/total_bits [23]),
	.I1(\top/processor/total_bits [22]),
	.I2(\top/processor/total_bits [21]),
	.F(\top/processor/n11417_15 )
);
defparam \top/processor/n11417_s10 .INIT=8'h80;
LUT3 \top/processor/n11416_s10  (
	.I0(\top/processor/total_bits [24]),
	.I1(\top/processor/n11420_15 ),
	.I2(\top/processor/n11417_15 ),
	.F(\top/processor/n11416_15 )
);
defparam \top/processor/n11416_s10 .INIT=8'h80;
LUT4 \top/processor/n11415_s10  (
	.I0(\top/processor/total_bits [25]),
	.I1(\top/processor/total_bits [24]),
	.I2(\top/processor/n11420_15 ),
	.I3(\top/processor/n11417_15 ),
	.F(\top/processor/n11415_15 )
);
defparam \top/processor/n11415_s10 .INIT=16'h8000;
LUT2 \top/processor/n11414_s10  (
	.I0(\top/processor/total_bits [26]),
	.I1(\top/processor/n11415_15 ),
	.F(\top/processor/n11414_15 )
);
defparam \top/processor/n11414_s10 .INIT=4'h8;
LUT2 \top/processor/n11412_s10  (
	.I0(\top/processor/total_bits [28]),
	.I1(\top/processor/total_bits [27]),
	.F(\top/processor/n11412_15 )
);
defparam \top/processor/n11412_s10 .INIT=4'h8;
LUT3 \top/processor/n11411_s10  (
	.I0(\top/processor/total_bits [29]),
	.I1(\top/processor/total_bits [28]),
	.I2(\top/processor/total_bits [27]),
	.F(\top/processor/n11411_15 )
);
defparam \top/processor/n11411_s10 .INIT=8'h80;
LUT4 \top/processor/n11410_s10  (
	.I0(\top/processor/n11410_19 ),
	.I1(\top/processor/total_bits [25]),
	.I2(\top/processor/total_bits [24]),
	.I3(\top/processor/n11420_15 ),
	.F(\top/processor/n11410_15 )
);
defparam \top/processor/n11410_s10 .INIT=16'h8000;
LUT2 \top/processor/n11409_s10  (
	.I0(\top/processor/total_bits [31]),
	.I1(\top/processor/n11410_15 ),
	.F(\top/processor/n11409_15 )
);
defparam \top/processor/n11409_s10 .INIT=4'h8;
LUT4 \top/processor/n11407_s10  (
	.I0(\top/processor/total_bits [33]),
	.I1(\top/processor/total_bits [32]),
	.I2(\top/processor/total_bits [31]),
	.I3(\top/processor/n11410_15 ),
	.F(\top/processor/n11407_15 )
);
defparam \top/processor/n11407_s10 .INIT=16'h8000;
LUT4 \top/processor/n11405_s10  (
	.I0(\top/processor/total_bits [35]),
	.I1(\top/processor/total_bits [25]),
	.I2(\top/processor/n11420_15 ),
	.I3(\top/processor/n11405_16 ),
	.F(\top/processor/n11405_15 )
);
defparam \top/processor/n11405_s10 .INIT=16'h8000;
LUT2 \top/processor/n11403_s10  (
	.I0(\top/processor/total_bits [37]),
	.I1(\top/processor/total_bits [36]),
	.F(\top/processor/n11403_15 )
);
defparam \top/processor/n11403_s10 .INIT=4'h8;
LUT4 \top/processor/n11400_s10  (
	.I0(\top/processor/total_bits [40]),
	.I1(\top/processor/total_bits [39]),
	.I2(\top/processor/total_bits [38]),
	.I3(\top/processor/n11403_15 ),
	.F(\top/processor/n11400_15 )
);
defparam \top/processor/n11400_s10 .INIT=16'h8000;
LUT3 \top/processor/n11399_s10  (
	.I0(\top/processor/total_bits [41]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/n11400_15 ),
	.F(\top/processor/n11399_15 )
);
defparam \top/processor/n11399_s10 .INIT=8'h80;
LUT4 \top/processor/n11398_s10  (
	.I0(\top/processor/total_bits [42]),
	.I1(\top/processor/total_bits [41]),
	.I2(\top/processor/n11405_15 ),
	.I3(\top/processor/n11400_15 ),
	.F(\top/processor/n11398_15 )
);
defparam \top/processor/n11398_s10 .INIT=16'h8000;
LUT4 \top/processor/n11396_s10  (
	.I0(\top/processor/total_bits [44]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/n11400_15 ),
	.I3(\top/processor/n11396_16 ),
	.F(\top/processor/n11396_15 )
);
defparam \top/processor/n11396_s10 .INIT=16'h8000;
LUT4 \top/processor/n11395_s10  (
	.I0(\top/processor/total_bits [45]),
	.I1(\top/processor/total_bits [44]),
	.I2(\top/processor/n11400_15 ),
	.I3(\top/processor/n11396_16 ),
	.F(\top/processor/n11395_15 )
);
defparam \top/processor/n11395_s10 .INIT=16'h8000;
LUT3 \top/processor/n11394_s10  (
	.I0(\top/processor/total_bits [46]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/n11395_15 ),
	.F(\top/processor/n11394_15 )
);
defparam \top/processor/n11394_s10 .INIT=8'h80;
LUT3 \top/processor/n11392_s10  (
	.I0(\top/processor/n11405_15 ),
	.I1(\top/processor/n11395_15 ),
	.I2(\top/processor/n11392_16 ),
	.F(\top/processor/n11392_15 )
);
defparam \top/processor/n11392_s10 .INIT=8'h80;
LUT2 \top/processor/n11390_s10  (
	.I0(\top/processor/n11405_15 ),
	.I1(\top/processor/n11390_16 ),
	.F(\top/processor/n11390_15 )
);
defparam \top/processor/n11390_s10 .INIT=4'h8;
LUT2 \top/processor/n11388_s10  (
	.I0(\top/processor/total_bits [52]),
	.I1(\top/processor/total_bits [51]),
	.F(\top/processor/n11388_15 )
);
defparam \top/processor/n11388_s10 .INIT=4'h8;
LUT4 \top/processor/n11387_s10  (
	.I0(\top/processor/total_bits [53]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/n11390_16 ),
	.I3(\top/processor/n11388_15 ),
	.F(\top/processor/n11387_15 )
);
defparam \top/processor/n11387_s10 .INIT=16'h8000;
LUT3 \top/processor/n11385_s10  (
	.I0(\top/processor/n11405_15 ),
	.I1(\top/processor/n11390_16 ),
	.I2(\top/processor/n11385_16 ),
	.F(\top/processor/n11385_15 )
);
defparam \top/processor/n11385_s10 .INIT=8'h80;
LUT2 \top/processor/n11383_s10  (
	.I0(\top/processor/total_bits [57]),
	.I1(\top/processor/total_bits [56]),
	.F(\top/processor/n11383_15 )
);
defparam \top/processor/n11383_s10 .INIT=4'h8;
LUT4 \top/processor/n11382_s10  (
	.I0(\top/processor/n11382_18 ),
	.I1(\top/processor/total_bits [58]),
	.I2(\top/processor/n11405_15 ),
	.I3(\top/processor/n11390_16 ),
	.F(\top/processor/n11382_15 )
);
defparam \top/processor/n11382_s10 .INIT=16'h8000;
LUT2 \top/processor/n11380_s10  (
	.I0(\top/processor/total_bits [60]),
	.I1(\top/processor/total_bits [59]),
	.F(\top/processor/n11380_15 )
);
defparam \top/processor/n11380_s10 .INIT=4'h8;
LUT2 \top/processor/n11377_s10  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/n11374_20 ),
	.F(\top/processor/n11377_15 )
);
defparam \top/processor/n11377_s10 .INIT=4'h1;
LUT4 \top/processor/n11376_s10  (
	.I0(\top/processor/n11374_20 ),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [1]),
	.I3(\top/processor/n11376_16 ),
	.F(\top/processor/n11376_15 )
);
defparam \top/processor/n11376_s10 .INIT=16'h00EB;
LUT3 \top/processor/n11375_s10  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/byte_index [2]),
	.F(\top/processor/n11375_15 )
);
defparam \top/processor/n11375_s10 .INIT=8'h78;
LUT4 \top/processor/n11375_s11  (
	.I0(\top/processor/pad_index [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/n11374_20 ),
	.I3(\top/processor/pad_index [2]),
	.F(\top/processor/n11375_16 )
);
defparam \top/processor/n11375_s11 .INIT=16'h0708;
LUT3 \top/processor/n11374_s12  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/block_buffer_391_9 ),
	.I2(\top/processor/n10817_15 ),
	.F(\top/processor/n11374_17 )
);
defparam \top/processor/n11374_s12 .INIT=8'h60;
LUT3 \top/processor/n11373_s10  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/block_buffer_391_9 ),
	.I2(\top/processor/byte_index [4]),
	.F(\top/processor/n11373_15 )
);
defparam \top/processor/n11373_s10 .INIT=8'h78;
LUT4 \top/processor/n11373_s11  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/block_buffer_455_9 ),
	.I2(\top/processor/n11374_20 ),
	.I3(\top/processor/pad_index [4]),
	.F(\top/processor/n11373_16 )
);
defparam \top/processor/n11373_s11 .INIT=16'h0708;
LUT4 \top/processor/n11372_s10  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [3]),
	.I2(\top/processor/block_buffer_391_9 ),
	.I3(\top/processor/byte_index [5]),
	.F(\top/processor/n11372_15 )
);
defparam \top/processor/n11372_s10 .INIT=16'h807F;
LUT4 \top/processor/n11372_s11  (
	.I0(\top/processor/need_length_block ),
	.I1(\top/processor/n11374_18 ),
	.I2(\top/processor/block_buffer_455_9 ),
	.I3(\top/processor/pad_index [5]),
	.F(\top/processor/n11372_16 )
);
defparam \top/processor/n11372_s11 .INIT=16'hC43F;
LUT2 \top/processor/n11370_s13  (
	.I0(\top/state_0 [1]),
	.I1(\top/state_0 [0]),
	.F(\top/processor/n11370_19 )
);
defparam \top/processor/n11370_s13 .INIT=4'h4;
LUT2 \top/processor/n11362_s12  (
	.I0(\top/processor/seen_last ),
	.I1(\top/processor/need_length_block ),
	.F(\top/processor/n11362_19 )
);
defparam \top/processor/n11362_s12 .INIT=4'h8;
LUT4 \top/processor/state_1_s6  (
	.I0(\top/processor/seen_last ),
	.I1(\top/data_last ),
	.I2(\top/state_0 [0]),
	.I3(\top/data_valid ),
	.F(\top/processor/state_1_10 )
);
defparam \top/processor/state_1_s6 .INIT=16'hC35C;
LUT3 \top/processor/block_buffer_511_s8  (
	.I0(\top/processor/block_buffer_503_9 ),
	.I1(\top/processor/block_buffer_319_15 ),
	.I2(\top/processor/n7631_8 ),
	.F(\top/processor/block_buffer_511_12 )
);
defparam \top/processor/block_buffer_511_s8 .INIT=8'h07;
LUT3 \top/processor/block_buffer_511_s9  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [3]),
	.I2(\top/processor/byte_index [5]),
	.F(\top/processor/block_buffer_511_13 )
);
defparam \top/processor/block_buffer_511_s9 .INIT=8'h01;
LUT4 \top/processor/block_buffer_447_s6  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [5]),
	.I2(\top/processor/byte_index [3]),
	.I3(\top/processor/block_buffer_319_9 ),
	.F(\top/processor/block_buffer_447_10 )
);
defparam \top/processor/block_buffer_447_s6 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_447_s7  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/block_buffer_447_10 ),
	.I2(\top/processor/block_buffer_63_10 ),
	.I3(\top/processor/block_buffer_447_12 ),
	.F(\top/processor/block_buffer_447_11 )
);
defparam \top/processor/block_buffer_447_s7 .INIT=16'hE000;
LUT4 \top/processor/block_buffer_439_s8  (
	.I0(\top/processor/pad_index [4]),
	.I1(\top/processor/pad_index [5]),
	.I2(\top/state_0 [1]),
	.I3(\top/processor/pad_index [3]),
	.F(\top/processor/block_buffer_439_12 )
);
defparam \top/processor/block_buffer_439_s8 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_423_s7  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [2]),
	.I2(\top/processor/pad_index [1]),
	.I3(\top/processor/pad_index [0]),
	.F(\top/processor/block_buffer_423_11 )
);
defparam \top/processor/block_buffer_423_s7 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_407_s7  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [1]),
	.I2(\top/processor/pad_index [0]),
	.I3(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_407_11 )
);
defparam \top/processor/block_buffer_407_s7 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_383_s6  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/byte_index [5]),
	.I2(\top/processor/byte_index [4]),
	.I3(\top/processor/block_buffer_319_9 ),
	.F(\top/processor/block_buffer_383_10 )
);
defparam \top/processor/block_buffer_383_s6 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_383_s7  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [5]),
	.I2(\top/state_0 [1]),
	.I3(\top/processor/block_buffer_319_15 ),
	.F(\top/processor/block_buffer_383_11 )
);
defparam \top/processor/block_buffer_383_s7 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_375_s7  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [5]),
	.I2(\top/processor/pad_index [4]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/block_buffer_375_11 )
);
defparam \top/processor/block_buffer_375_s7 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_255_s6  (
	.I0(\top/processor/byte_index [4]),
	.I1(\top/processor/byte_index [3]),
	.I2(\top/processor/byte_index [5]),
	.I3(\top/processor/block_buffer_319_9 ),
	.F(\top/processor/block_buffer_255_10 )
);
defparam \top/processor/block_buffer_255_s6 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_255_s7  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [4]),
	.I2(\top/state_0 [1]),
	.I3(\top/processor/block_buffer_319_15 ),
	.F(\top/processor/block_buffer_255_11 )
);
defparam \top/processor/block_buffer_255_s7 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_247_s7  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [4]),
	.I2(\top/state_0 [1]),
	.I3(\top/processor/pad_index [5]),
	.F(\top/processor/block_buffer_247_11 )
);
defparam \top/processor/block_buffer_247_s7 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_191_s7  (
	.I0(\top/processor/pad_index [4]),
	.I1(\top/processor/pad_index [3]),
	.I2(\top/state_0 [1]),
	.I3(\top/processor/pad_index [5]),
	.F(\top/processor/block_buffer_191_11 )
);
defparam \top/processor/block_buffer_191_s7 .INIT=16'h4000;
LUT4 \top/processor/block_buffer_127_s7  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/pad_index [4]),
	.I3(\top/processor/pad_index [5]),
	.F(\top/processor/block_buffer_127_11 )
);
defparam \top/processor/block_buffer_127_s7 .INIT=16'h4000;
LUT4 \top/processor/n11420_s11  (
	.I0(\top/processor/total_bits [18]),
	.I1(\top/processor/total_bits [17]),
	.I2(\top/processor/total_bits [16]),
	.I3(\top/processor/n11425_15 ),
	.F(\top/processor/n11420_16 )
);
defparam \top/processor/n11420_s11 .INIT=16'h8000;
LUT4 \top/processor/n11405_s11  (
	.I0(\top/processor/n11405_17 ),
	.I1(\top/processor/total_bits [34]),
	.I2(\top/processor/total_bits [33]),
	.I3(\top/processor/n11410_17 ),
	.F(\top/processor/n11405_16 )
);
defparam \top/processor/n11405_s11 .INIT=16'h8000;
LUT3 \top/processor/n11396_s11  (
	.I0(\top/processor/total_bits [43]),
	.I1(\top/processor/total_bits [42]),
	.I2(\top/processor/total_bits [41]),
	.F(\top/processor/n11396_16 )
);
defparam \top/processor/n11396_s11 .INIT=8'h80;
LUT3 \top/processor/n11392_s11  (
	.I0(\top/processor/total_bits [48]),
	.I1(\top/processor/total_bits [47]),
	.I2(\top/processor/total_bits [46]),
	.F(\top/processor/n11392_16 )
);
defparam \top/processor/n11392_s11 .INIT=8'h80;
LUT4 \top/processor/n11390_s11  (
	.I0(\top/processor/total_bits [50]),
	.I1(\top/processor/total_bits [49]),
	.I2(\top/processor/n11395_15 ),
	.I3(\top/processor/n11392_16 ),
	.F(\top/processor/n11390_16 )
);
defparam \top/processor/n11390_s11 .INIT=16'h8000;
LUT4 \top/processor/n11385_s11  (
	.I0(\top/processor/total_bits [55]),
	.I1(\top/processor/total_bits [54]),
	.I2(\top/processor/total_bits [53]),
	.I3(\top/processor/n11388_15 ),
	.F(\top/processor/n11385_16 )
);
defparam \top/processor/n11385_s11 .INIT=16'h8000;
LUT3 \top/processor/n11376_s11  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/processor/n10817_15 ),
	.F(\top/processor/n11376_16 )
);
defparam \top/processor/n11376_s11 .INIT=8'h60;
LUT2 \top/processor/n11374_s13  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [4]),
	.F(\top/processor/n11374_18 )
);
defparam \top/processor/n11374_s13 .INIT=4'h8;
LUT4 \top/processor/block_buffer_447_s8  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [4]),
	.I2(\top/processor/pad_index [5]),
	.I3(\top/state_0 [1]),
	.F(\top/processor/block_buffer_447_12 )
);
defparam \top/processor/block_buffer_447_s8 .INIT=16'h0100;
LUT4 \top/processor/n11410_s12  (
	.I0(\top/processor/total_bits [30]),
	.I1(\top/processor/total_bits [29]),
	.I2(\top/processor/total_bits [26]),
	.I3(\top/processor/n11412_15 ),
	.F(\top/processor/n11410_17 )
);
defparam \top/processor/n11410_s12 .INIT=16'h8000;
LUT4 \top/processor/n11405_s12  (
	.I0(\top/processor/total_bits [32]),
	.I1(\top/processor/total_bits [31]),
	.I2(\top/processor/total_bits [24]),
	.I3(\top/processor/n11417_15 ),
	.F(\top/processor/n11405_17 )
);
defparam \top/processor/n11405_s12 .INIT=16'h8000;
LUT3 \top/processor/n11379_s11  (
	.I0(\top/processor/total_bits [61]),
	.I1(\top/processor/total_bits [60]),
	.I2(\top/processor/total_bits [59]),
	.F(\top/processor/n11379_17 )
);
defparam \top/processor/n11379_s11 .INIT=8'h80;
LUT3 \top/processor/n11382_s12  (
	.I0(\top/processor/n11385_16 ),
	.I1(\top/processor/total_bits [57]),
	.I2(\top/processor/total_bits [56]),
	.F(\top/processor/n11382_18 )
);
defparam \top/processor/n11382_s12 .INIT=8'h80;
LUT4 \top/processor/n11409_s11  (
	.I0(\top/processor/total_bits [32]),
	.I1(\top/processor/total_bits [31]),
	.I2(\top/processor/n11410_15 ),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11409_17 )
);
defparam \top/processor/n11409_s11 .INIT=16'h6A00;
LUT4 \top/processor/n9790_s7  (
	.I0(\top/processor/n9790_11 ),
	.I1(\top/state_0 [2]),
	.I2(\top/processor/core_busy ),
	.I3(\top/processor/block_ready ),
	.F(\top/processor/n9790_13 )
);
defparam \top/processor/n9790_s7 .INIT=16'h0200;
LUT4 \top/processor/block_buffer_399_s8  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [1]),
	.I3(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_399_13 )
);
defparam \top/processor/block_buffer_399_s8 .INIT=16'h1000;
LUT4 \top/processor/block_buffer_431_s8  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [2]),
	.I3(\top/processor/pad_index [1]),
	.F(\top/processor/block_buffer_431_13 )
);
defparam \top/processor/block_buffer_431_s8 .INIT=16'h0100;
LUT4 \top/processor/n11390_s12  (
	.I0(\top/processor/total_bits [51]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/n11390_16 ),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11390_18 )
);
defparam \top/processor/n11390_s12 .INIT=16'h6A00;
LUT4 \top/processor/n11402_s11  (
	.I0(\top/processor/total_bits [38]),
	.I1(\top/processor/n11405_15 ),
	.I2(\top/processor/total_bits [37]),
	.I3(\top/processor/total_bits [36]),
	.F(\top/processor/n11402_17 )
);
defparam \top/processor/n11402_s11 .INIT=16'h8000;
LUT4 \top/processor/n11427_s11  (
	.I0(\top/processor/total_bits [13]),
	.I1(\top/processor/n11430_15 ),
	.I2(\top/processor/total_bits [12]),
	.I3(\top/processor/total_bits [11]),
	.F(\top/processor/n11427_17 )
);
defparam \top/processor/n11427_s11 .INIT=16'h8000;
LUT4 \top/processor/block_buffer_319_s10  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [1]),
	.I3(\top/processor/pad_index [2]),
	.F(\top/processor/block_buffer_319_15 )
);
defparam \top/processor/block_buffer_319_s10 .INIT=16'h0001;
LUT4 \top/processor/block_buffer_263_s7  (
	.I0(\top/state_0 [0]),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/pad_index [3]),
	.I3(\top/processor/pad_index [4]),
	.F(\top/processor/block_buffer_263_12 )
);
defparam \top/processor/block_buffer_263_s7 .INIT=16'h4000;
LUT4 \top/processor/block_buffer_319_s11  (
	.I0(\top/processor/pad_index [5]),
	.I1(\top/state_0 [1]),
	.I2(\top/processor/pad_index [3]),
	.I3(\top/processor/pad_index [4]),
	.F(\top/processor/block_buffer_319_17 )
);
defparam \top/processor/block_buffer_319_s11 .INIT=16'h4000;
LUT4 \top/processor/n11374_s14  (
	.I0(\top/processor/need_length_block ),
	.I1(\top/processor/pad_index [5]),
	.I2(\top/processor/pad_index [3]),
	.I3(\top/processor/pad_index [4]),
	.F(\top/processor/n11374_20 )
);
defparam \top/processor/n11374_s14 .INIT=16'h4000;
LUT4 \top/processor/n11414_s11  (
	.I0(\top/processor/total_bits [27]),
	.I1(\top/processor/total_bits [26]),
	.I2(\top/processor/n11415_15 ),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11414_17 )
);
defparam \top/processor/n11414_s11 .INIT=16'h6A00;
LUT4 \top/processor/n11410_s13  (
	.I0(\top/processor/total_bits [23]),
	.I1(\top/processor/total_bits [22]),
	.I2(\top/processor/total_bits [21]),
	.I3(\top/processor/n11410_17 ),
	.F(\top/processor/n11410_19 )
);
defparam \top/processor/n11410_s13 .INIT=16'h8000;
LUT4 \top/processor/core_busy_s3  (
	.I0(\top/processor/core_ready_prev ),
	.I1(\top/processor/core_ready ),
	.I2(\top/processor/n9790_15 ),
	.I3(\top/processor/n9790_13 ),
	.F(\top/processor/core_busy_8 )
);
defparam \top/processor/core_busy_s3 .INIT=16'hFF40;
LUT3 \top/processor/n9790_s8  (
	.I0(\top/state_0 [2]),
	.I1(\top/state_0 [0]),
	.I2(\top/state_0 [1]),
	.F(\top/processor/n9790_15 )
);
defparam \top/processor/n9790_s8 .INIT=8'h40;
LUT4 \top/processor/n11424_s11  (
	.I0(\top/processor/total_bits [16]),
	.I1(\top/processor/total_bits [10]),
	.I2(\top/processor/n11431_15 ),
	.I3(\top/processor/n11425_15 ),
	.F(\top/processor/n11424_17 )
);
defparam \top/processor/n11424_s11 .INIT=16'h8000;
LUT4 \top/processor/n11430_s11  (
	.I0(\top/processor/total_bits [11]),
	.I1(\top/processor/total_bits [10]),
	.I2(\top/processor/n11431_15 ),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11430_17 )
);
defparam \top/processor/n11430_s11 .INIT=16'h6A00;
LUT3 \top/processor/n7631_s4  (
	.I0(\top/data_valid ),
	.I1(\top/state_0 [1]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n7631_8 )
);
defparam \top/processor/n7631_s4 .INIT=8'h20;
LUT3 \top/processor/n11365_s12  (
	.I0(\top/state_0 [1]),
	.I1(\top/state_0 [0]),
	.I2(\top/processor/n11372_15 ),
	.F(\top/processor/n11365_19 )
);
defparam \top/processor/n11365_s12 .INIT=8'h04;
LUT4 \top/processor/n11367_s12  (
	.I0(\top/processor/byte_index [3]),
	.I1(\top/processor/block_buffer_391_9 ),
	.I2(\top/state_0 [1]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11367_19 )
);
defparam \top/processor/n11367_s12 .INIT=16'h0600;
LUT4 \top/processor/n11369_s12  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/processor/byte_index [1]),
	.I2(\top/state_0 [1]),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11369_19 )
);
defparam \top/processor/n11369_s12 .INIT=16'h0600;
LUT3 \top/processor/n11370_s14  (
	.I0(\top/processor/byte_index [0]),
	.I1(\top/state_0 [1]),
	.I2(\top/state_0 [0]),
	.F(\top/processor/n11370_21 )
);
defparam \top/processor/n11370_s14 .INIT=8'h10;
LUT4 \top/processor/n7631_s5  (
	.I0(\top/processor/pad_index [5]),
	.I1(\top/processor/block_buffer_263_12 ),
	.I2(\top/processor/need_length_block ),
	.I3(\top/processor/block_buffer_511_9 ),
	.F(\top/processor/n7631_10 )
);
defparam \top/processor/n7631_s5 .INIT=16'h00F7;
LUT4 \top/processor/n7631_s6  (
	.I0(\top/processor/block_buffer_391_9 ),
	.I1(\top/processor/byte_index [4]),
	.I2(\top/processor/byte_index [3]),
	.I3(\top/processor/byte_index [5]),
	.F(\top/processor/n7631_12 )
);
defparam \top/processor/n7631_s6 .INIT=16'h8000;
LUT4 \top/processor/n11374_s15  (
	.I0(\top/processor/pad_index [3]),
	.I1(\top/processor/pad_index [0]),
	.I2(\top/processor/pad_index [1]),
	.I3(\top/processor/pad_index [2]),
	.F(\top/processor/n11374_22 )
);
defparam \top/processor/n11374_s15 .INIT=16'h6AAA;
LUT3 \top/processor/block_buffer_495_s8  (
	.I0(\top/state_0 [0]),
	.I1(\top/processor/n11374_20 ),
	.I2(\top/processor/block_buffer_503_9 ),
	.F(\top/processor/block_buffer_495_13 )
);
defparam \top/processor/block_buffer_495_s8 .INIT=8'h10;
LUT4 \top/processor/block_buffer_7_s6  (
	.I0(\top/processor/n7631_10 ),
	.I1(\top/processor/block_buffer_7_9 ),
	.I2(\top/state_0 [2]),
	.I3(rst),
	.F(\top/processor/block_buffer_7_11 )
);
defparam \top/processor/block_buffer_7_s6 .INIT=16'h0007;
LUT4 \top/processor/block_buffer_255_s8  (
	.I0(\top/processor/block_buffer_511_9 ),
	.I1(\top/processor/block_buffer_255_9 ),
	.I2(\top/state_0 [2]),
	.I3(rst),
	.F(\top/processor/block_buffer_255_13 )
);
defparam \top/processor/block_buffer_255_s8 .INIT=16'h000E;
LUT4 \top/processor/block_buffer_383_s8  (
	.I0(\top/processor/block_buffer_511_9 ),
	.I1(\top/processor/block_buffer_383_9 ),
	.I2(\top/state_0 [2]),
	.I3(rst),
	.F(\top/processor/block_buffer_383_13 )
);
defparam \top/processor/block_buffer_383_s8 .INIT=16'h000E;
LUT3 \top/processor/block_buffer_447_s9  (
	.I0(\top/processor/block_buffer_447_9 ),
	.I1(\top/state_0 [2]),
	.I2(rst),
	.F(\top/processor/block_buffer_447_14 )
);
defparam \top/processor/block_buffer_447_s9 .INIT=8'h01;
LUT4 \top/processor/block_buffer_511_s10  (
	.I0(\top/processor/block_buffer_511_9 ),
	.I1(\top/processor/block_buffer_511_10 ),
	.I2(\top/state_0 [2]),
	.I3(rst),
	.F(\top/processor/block_buffer_511_15 )
);
defparam \top/processor/block_buffer_511_s10 .INIT=16'h000E;
LUT4 \top/processor/n11378_s11  (
	.I0(\top/processor/total_bits [62]),
	.I1(\top/processor/total_bits [61]),
	.I2(\top/processor/total_bits [60]),
	.I3(\top/processor/total_bits [59]),
	.F(\top/processor/n11378_17 )
);
defparam \top/processor/n11378_s11 .INIT=16'h8000;
LUT4 \top/processor/n11421_s11  (
	.I0(\top/processor/total_bits [19]),
	.I1(\top/processor/total_bits [18]),
	.I2(\top/processor/total_bits [17]),
	.I3(\top/processor/n11424_17 ),
	.F(\top/processor/n11421_17 )
);
defparam \top/processor/n11421_s11 .INIT=16'h8000;
LUT4 \top/processor/n11423_s11  (
	.I0(\top/processor/total_bits [18]),
	.I1(\top/processor/total_bits [17]),
	.I2(\top/processor/n11424_17 ),
	.I3(\top/state_0 [0]),
	.F(\top/processor/n11423_17 )
);
defparam \top/processor/n11423_s11 .INIT=16'h6A00;
DFFCE \top/processor/state_1_s0  (
	.D(\top/processor/n11363_16 ),
	.CLK(clk),
	.CE(\top/processor/state_0_10 ),
	.CLEAR(rst),
	.Q(\top/state_0 [1])
);
defparam \top/processor/state_1_s0 .INIT=1'b0;
DFFCE \top/processor/state_0_s0  (
	.D(\top/processor/n11364_27 ),
	.CLK(clk),
	.CE(\top/processor/state_0_10 ),
	.CLEAR(rst),
	.Q(\top/state_0 [0])
);
defparam \top/processor/state_0_s0 .INIT=1'b0;
DFFCE \top/processor/byte_index_5_s0  (
	.D(\top/processor/n11365_19 ),
	.CLK(clk),
	.CE(\top/processor/byte_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/byte_index [5])
);
defparam \top/processor/byte_index_5_s0 .INIT=1'b0;
DFFCE \top/processor/byte_index_4_s0  (
	.D(\top/processor/n11366_17 ),
	.CLK(clk),
	.CE(\top/processor/byte_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/byte_index [4])
);
defparam \top/processor/byte_index_4_s0 .INIT=1'b0;
DFFCE \top/processor/byte_index_3_s0  (
	.D(\top/processor/n11367_19 ),
	.CLK(clk),
	.CE(\top/processor/byte_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/byte_index [3])
);
defparam \top/processor/byte_index_3_s0 .INIT=1'b0;
DFFCE \top/processor/byte_index_2_s0  (
	.D(\top/processor/n11368_17 ),
	.CLK(clk),
	.CE(\top/processor/byte_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/byte_index [2])
);
defparam \top/processor/byte_index_2_s0 .INIT=1'b0;
DFFCE \top/processor/byte_index_1_s0  (
	.D(\top/processor/n11369_19 ),
	.CLK(clk),
	.CE(\top/processor/byte_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/byte_index [1])
);
defparam \top/processor/byte_index_1_s0 .INIT=1'b0;
DFFCE \top/processor/byte_index_0_s0  (
	.D(\top/processor/n11370_21 ),
	.CLK(clk),
	.CE(\top/processor/byte_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/byte_index [0])
);
defparam \top/processor/byte_index_0_s0 .INIT=1'b0;
DFFCE \top/processor/block_ready_s0  (
	.D(\top/processor/n7631_3 ),
	.CLK(clk),
	.CE(\top/processor/block_ready_8 ),
	.CLEAR(rst),
	.Q(\top/processor/block_ready )
);
defparam \top/processor/block_ready_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_511_s0  (
	.D(\top/processor/block_buffer [511]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [511])
);
defparam \top/processor/core_block_511_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_510_s0  (
	.D(\top/processor/block_buffer [510]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [510])
);
defparam \top/processor/core_block_510_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_509_s0  (
	.D(\top/processor/block_buffer [509]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [509])
);
defparam \top/processor/core_block_509_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_508_s0  (
	.D(\top/processor/block_buffer [508]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [508])
);
defparam \top/processor/core_block_508_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_507_s0  (
	.D(\top/processor/block_buffer [507]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [507])
);
defparam \top/processor/core_block_507_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_506_s0  (
	.D(\top/processor/block_buffer [506]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [506])
);
defparam \top/processor/core_block_506_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_505_s0  (
	.D(\top/processor/block_buffer [505]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [505])
);
defparam \top/processor/core_block_505_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_504_s0  (
	.D(\top/processor/block_buffer [504]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [504])
);
defparam \top/processor/core_block_504_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_503_s0  (
	.D(\top/processor/block_buffer [503]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [503])
);
defparam \top/processor/core_block_503_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_502_s0  (
	.D(\top/processor/block_buffer [502]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [502])
);
defparam \top/processor/core_block_502_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_501_s0  (
	.D(\top/processor/block_buffer [501]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [501])
);
defparam \top/processor/core_block_501_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_500_s0  (
	.D(\top/processor/block_buffer [500]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [500])
);
defparam \top/processor/core_block_500_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_499_s0  (
	.D(\top/processor/block_buffer [499]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [499])
);
defparam \top/processor/core_block_499_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_498_s0  (
	.D(\top/processor/block_buffer [498]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [498])
);
defparam \top/processor/core_block_498_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_497_s0  (
	.D(\top/processor/block_buffer [497]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [497])
);
defparam \top/processor/core_block_497_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_496_s0  (
	.D(\top/processor/block_buffer [496]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [496])
);
defparam \top/processor/core_block_496_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_495_s0  (
	.D(\top/processor/block_buffer [495]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [495])
);
defparam \top/processor/core_block_495_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_494_s0  (
	.D(\top/processor/block_buffer [494]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [494])
);
defparam \top/processor/core_block_494_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_493_s0  (
	.D(\top/processor/block_buffer [493]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [493])
);
defparam \top/processor/core_block_493_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_492_s0  (
	.D(\top/processor/block_buffer [492]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [492])
);
defparam \top/processor/core_block_492_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_491_s0  (
	.D(\top/processor/block_buffer [491]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [491])
);
defparam \top/processor/core_block_491_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_490_s0  (
	.D(\top/processor/block_buffer [490]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [490])
);
defparam \top/processor/core_block_490_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_489_s0  (
	.D(\top/processor/block_buffer [489]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [489])
);
defparam \top/processor/core_block_489_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_488_s0  (
	.D(\top/processor/block_buffer [488]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [488])
);
defparam \top/processor/core_block_488_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_487_s0  (
	.D(\top/processor/block_buffer [487]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [487])
);
defparam \top/processor/core_block_487_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_486_s0  (
	.D(\top/processor/block_buffer [486]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [486])
);
defparam \top/processor/core_block_486_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_485_s0  (
	.D(\top/processor/block_buffer [485]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [485])
);
defparam \top/processor/core_block_485_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_484_s0  (
	.D(\top/processor/block_buffer [484]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [484])
);
defparam \top/processor/core_block_484_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_483_s0  (
	.D(\top/processor/block_buffer [483]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [483])
);
defparam \top/processor/core_block_483_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_482_s0  (
	.D(\top/processor/block_buffer [482]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [482])
);
defparam \top/processor/core_block_482_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_481_s0  (
	.D(\top/processor/block_buffer [481]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [481])
);
defparam \top/processor/core_block_481_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_480_s0  (
	.D(\top/processor/block_buffer [480]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [480])
);
defparam \top/processor/core_block_480_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_479_s0  (
	.D(\top/processor/block_buffer [479]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [479])
);
defparam \top/processor/core_block_479_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_478_s0  (
	.D(\top/processor/block_buffer [478]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [478])
);
defparam \top/processor/core_block_478_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_477_s0  (
	.D(\top/processor/block_buffer [477]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [477])
);
defparam \top/processor/core_block_477_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_476_s0  (
	.D(\top/processor/block_buffer [476]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [476])
);
defparam \top/processor/core_block_476_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_475_s0  (
	.D(\top/processor/block_buffer [475]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [475])
);
defparam \top/processor/core_block_475_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_474_s0  (
	.D(\top/processor/block_buffer [474]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [474])
);
defparam \top/processor/core_block_474_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_473_s0  (
	.D(\top/processor/block_buffer [473]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [473])
);
defparam \top/processor/core_block_473_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_472_s0  (
	.D(\top/processor/block_buffer [472]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [472])
);
defparam \top/processor/core_block_472_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_471_s0  (
	.D(\top/processor/block_buffer [471]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [471])
);
defparam \top/processor/core_block_471_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_470_s0  (
	.D(\top/processor/block_buffer [470]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [470])
);
defparam \top/processor/core_block_470_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_469_s0  (
	.D(\top/processor/block_buffer [469]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [469])
);
defparam \top/processor/core_block_469_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_468_s0  (
	.D(\top/processor/block_buffer [468]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [468])
);
defparam \top/processor/core_block_468_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_467_s0  (
	.D(\top/processor/block_buffer [467]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [467])
);
defparam \top/processor/core_block_467_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_466_s0  (
	.D(\top/processor/block_buffer [466]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [466])
);
defparam \top/processor/core_block_466_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_465_s0  (
	.D(\top/processor/block_buffer [465]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [465])
);
defparam \top/processor/core_block_465_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_464_s0  (
	.D(\top/processor/block_buffer [464]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [464])
);
defparam \top/processor/core_block_464_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_463_s0  (
	.D(\top/processor/block_buffer [463]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [463])
);
defparam \top/processor/core_block_463_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_462_s0  (
	.D(\top/processor/block_buffer [462]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [462])
);
defparam \top/processor/core_block_462_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_461_s0  (
	.D(\top/processor/block_buffer [461]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [461])
);
defparam \top/processor/core_block_461_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_460_s0  (
	.D(\top/processor/block_buffer [460]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [460])
);
defparam \top/processor/core_block_460_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_459_s0  (
	.D(\top/processor/block_buffer [459]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [459])
);
defparam \top/processor/core_block_459_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_458_s0  (
	.D(\top/processor/block_buffer [458]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [458])
);
defparam \top/processor/core_block_458_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_457_s0  (
	.D(\top/processor/block_buffer [457]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [457])
);
defparam \top/processor/core_block_457_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_456_s0  (
	.D(\top/processor/block_buffer [456]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [456])
);
defparam \top/processor/core_block_456_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_455_s0  (
	.D(\top/processor/block_buffer [455]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [455])
);
defparam \top/processor/core_block_455_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_454_s0  (
	.D(\top/processor/block_buffer [454]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [454])
);
defparam \top/processor/core_block_454_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_453_s0  (
	.D(\top/processor/block_buffer [453]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [453])
);
defparam \top/processor/core_block_453_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_452_s0  (
	.D(\top/processor/block_buffer [452]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [452])
);
defparam \top/processor/core_block_452_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_451_s0  (
	.D(\top/processor/block_buffer [451]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [451])
);
defparam \top/processor/core_block_451_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_450_s0  (
	.D(\top/processor/block_buffer [450]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [450])
);
defparam \top/processor/core_block_450_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_449_s0  (
	.D(\top/processor/block_buffer [449]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [449])
);
defparam \top/processor/core_block_449_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_448_s0  (
	.D(\top/processor/block_buffer [448]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [448])
);
defparam \top/processor/core_block_448_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_447_s0  (
	.D(\top/processor/block_buffer [447]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [447])
);
defparam \top/processor/core_block_447_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_446_s0  (
	.D(\top/processor/block_buffer [446]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [446])
);
defparam \top/processor/core_block_446_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_445_s0  (
	.D(\top/processor/block_buffer [445]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [445])
);
defparam \top/processor/core_block_445_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_444_s0  (
	.D(\top/processor/block_buffer [444]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [444])
);
defparam \top/processor/core_block_444_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_443_s0  (
	.D(\top/processor/block_buffer [443]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [443])
);
defparam \top/processor/core_block_443_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_442_s0  (
	.D(\top/processor/block_buffer [442]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [442])
);
defparam \top/processor/core_block_442_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_441_s0  (
	.D(\top/processor/block_buffer [441]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [441])
);
defparam \top/processor/core_block_441_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_440_s0  (
	.D(\top/processor/block_buffer [440]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [440])
);
defparam \top/processor/core_block_440_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_439_s0  (
	.D(\top/processor/block_buffer [439]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [439])
);
defparam \top/processor/core_block_439_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_438_s0  (
	.D(\top/processor/block_buffer [438]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [438])
);
defparam \top/processor/core_block_438_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_437_s0  (
	.D(\top/processor/block_buffer [437]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [437])
);
defparam \top/processor/core_block_437_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_436_s0  (
	.D(\top/processor/block_buffer [436]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [436])
);
defparam \top/processor/core_block_436_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_435_s0  (
	.D(\top/processor/block_buffer [435]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [435])
);
defparam \top/processor/core_block_435_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_434_s0  (
	.D(\top/processor/block_buffer [434]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [434])
);
defparam \top/processor/core_block_434_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_433_s0  (
	.D(\top/processor/block_buffer [433]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [433])
);
defparam \top/processor/core_block_433_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_432_s0  (
	.D(\top/processor/block_buffer [432]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [432])
);
defparam \top/processor/core_block_432_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_431_s0  (
	.D(\top/processor/block_buffer [431]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [431])
);
defparam \top/processor/core_block_431_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_430_s0  (
	.D(\top/processor/block_buffer [430]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [430])
);
defparam \top/processor/core_block_430_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_429_s0  (
	.D(\top/processor/block_buffer [429]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [429])
);
defparam \top/processor/core_block_429_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_428_s0  (
	.D(\top/processor/block_buffer [428]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [428])
);
defparam \top/processor/core_block_428_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_427_s0  (
	.D(\top/processor/block_buffer [427]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [427])
);
defparam \top/processor/core_block_427_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_426_s0  (
	.D(\top/processor/block_buffer [426]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [426])
);
defparam \top/processor/core_block_426_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_425_s0  (
	.D(\top/processor/block_buffer [425]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [425])
);
defparam \top/processor/core_block_425_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_424_s0  (
	.D(\top/processor/block_buffer [424]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [424])
);
defparam \top/processor/core_block_424_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_423_s0  (
	.D(\top/processor/block_buffer [423]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [423])
);
defparam \top/processor/core_block_423_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_422_s0  (
	.D(\top/processor/block_buffer [422]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [422])
);
defparam \top/processor/core_block_422_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_421_s0  (
	.D(\top/processor/block_buffer [421]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [421])
);
defparam \top/processor/core_block_421_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_420_s0  (
	.D(\top/processor/block_buffer [420]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [420])
);
defparam \top/processor/core_block_420_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_419_s0  (
	.D(\top/processor/block_buffer [419]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [419])
);
defparam \top/processor/core_block_419_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_418_s0  (
	.D(\top/processor/block_buffer [418]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [418])
);
defparam \top/processor/core_block_418_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_417_s0  (
	.D(\top/processor/block_buffer [417]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [417])
);
defparam \top/processor/core_block_417_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_416_s0  (
	.D(\top/processor/block_buffer [416]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [416])
);
defparam \top/processor/core_block_416_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_415_s0  (
	.D(\top/processor/block_buffer [415]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [415])
);
defparam \top/processor/core_block_415_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_414_s0  (
	.D(\top/processor/block_buffer [414]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [414])
);
defparam \top/processor/core_block_414_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_413_s0  (
	.D(\top/processor/block_buffer [413]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [413])
);
defparam \top/processor/core_block_413_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_412_s0  (
	.D(\top/processor/block_buffer [412]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [412])
);
defparam \top/processor/core_block_412_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_411_s0  (
	.D(\top/processor/block_buffer [411]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [411])
);
defparam \top/processor/core_block_411_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_410_s0  (
	.D(\top/processor/block_buffer [410]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [410])
);
defparam \top/processor/core_block_410_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_409_s0  (
	.D(\top/processor/block_buffer [409]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [409])
);
defparam \top/processor/core_block_409_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_408_s0  (
	.D(\top/processor/block_buffer [408]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [408])
);
defparam \top/processor/core_block_408_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_407_s0  (
	.D(\top/processor/block_buffer [407]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [407])
);
defparam \top/processor/core_block_407_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_406_s0  (
	.D(\top/processor/block_buffer [406]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [406])
);
defparam \top/processor/core_block_406_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_405_s0  (
	.D(\top/processor/block_buffer [405]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [405])
);
defparam \top/processor/core_block_405_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_404_s0  (
	.D(\top/processor/block_buffer [404]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [404])
);
defparam \top/processor/core_block_404_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_403_s0  (
	.D(\top/processor/block_buffer [403]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [403])
);
defparam \top/processor/core_block_403_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_402_s0  (
	.D(\top/processor/block_buffer [402]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [402])
);
defparam \top/processor/core_block_402_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_401_s0  (
	.D(\top/processor/block_buffer [401]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [401])
);
defparam \top/processor/core_block_401_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_400_s0  (
	.D(\top/processor/block_buffer [400]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [400])
);
defparam \top/processor/core_block_400_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_399_s0  (
	.D(\top/processor/block_buffer [399]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [399])
);
defparam \top/processor/core_block_399_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_398_s0  (
	.D(\top/processor/block_buffer [398]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [398])
);
defparam \top/processor/core_block_398_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_397_s0  (
	.D(\top/processor/block_buffer [397]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [397])
);
defparam \top/processor/core_block_397_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_396_s0  (
	.D(\top/processor/block_buffer [396]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [396])
);
defparam \top/processor/core_block_396_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_395_s0  (
	.D(\top/processor/block_buffer [395]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [395])
);
defparam \top/processor/core_block_395_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_394_s0  (
	.D(\top/processor/block_buffer [394]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [394])
);
defparam \top/processor/core_block_394_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_393_s0  (
	.D(\top/processor/block_buffer [393]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [393])
);
defparam \top/processor/core_block_393_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_392_s0  (
	.D(\top/processor/block_buffer [392]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [392])
);
defparam \top/processor/core_block_392_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_391_s0  (
	.D(\top/processor/block_buffer [391]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [391])
);
defparam \top/processor/core_block_391_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_390_s0  (
	.D(\top/processor/block_buffer [390]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [390])
);
defparam \top/processor/core_block_390_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_389_s0  (
	.D(\top/processor/block_buffer [389]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [389])
);
defparam \top/processor/core_block_389_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_388_s0  (
	.D(\top/processor/block_buffer [388]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [388])
);
defparam \top/processor/core_block_388_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_387_s0  (
	.D(\top/processor/block_buffer [387]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [387])
);
defparam \top/processor/core_block_387_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_386_s0  (
	.D(\top/processor/block_buffer [386]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [386])
);
defparam \top/processor/core_block_386_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_385_s0  (
	.D(\top/processor/block_buffer [385]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [385])
);
defparam \top/processor/core_block_385_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_384_s0  (
	.D(\top/processor/block_buffer [384]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [384])
);
defparam \top/processor/core_block_384_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_383_s0  (
	.D(\top/processor/block_buffer [383]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [383])
);
defparam \top/processor/core_block_383_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_382_s0  (
	.D(\top/processor/block_buffer [382]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [382])
);
defparam \top/processor/core_block_382_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_381_s0  (
	.D(\top/processor/block_buffer [381]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [381])
);
defparam \top/processor/core_block_381_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_380_s0  (
	.D(\top/processor/block_buffer [380]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [380])
);
defparam \top/processor/core_block_380_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_379_s0  (
	.D(\top/processor/block_buffer [379]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [379])
);
defparam \top/processor/core_block_379_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_378_s0  (
	.D(\top/processor/block_buffer [378]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [378])
);
defparam \top/processor/core_block_378_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_377_s0  (
	.D(\top/processor/block_buffer [377]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [377])
);
defparam \top/processor/core_block_377_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_376_s0  (
	.D(\top/processor/block_buffer [376]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [376])
);
defparam \top/processor/core_block_376_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_375_s0  (
	.D(\top/processor/block_buffer [375]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [375])
);
defparam \top/processor/core_block_375_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_374_s0  (
	.D(\top/processor/block_buffer [374]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [374])
);
defparam \top/processor/core_block_374_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_373_s0  (
	.D(\top/processor/block_buffer [373]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [373])
);
defparam \top/processor/core_block_373_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_372_s0  (
	.D(\top/processor/block_buffer [372]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [372])
);
defparam \top/processor/core_block_372_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_371_s0  (
	.D(\top/processor/block_buffer [371]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [371])
);
defparam \top/processor/core_block_371_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_370_s0  (
	.D(\top/processor/block_buffer [370]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [370])
);
defparam \top/processor/core_block_370_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_369_s0  (
	.D(\top/processor/block_buffer [369]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [369])
);
defparam \top/processor/core_block_369_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_368_s0  (
	.D(\top/processor/block_buffer [368]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [368])
);
defparam \top/processor/core_block_368_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_367_s0  (
	.D(\top/processor/block_buffer [367]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [367])
);
defparam \top/processor/core_block_367_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_366_s0  (
	.D(\top/processor/block_buffer [366]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [366])
);
defparam \top/processor/core_block_366_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_365_s0  (
	.D(\top/processor/block_buffer [365]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [365])
);
defparam \top/processor/core_block_365_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_364_s0  (
	.D(\top/processor/block_buffer [364]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [364])
);
defparam \top/processor/core_block_364_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_363_s0  (
	.D(\top/processor/block_buffer [363]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [363])
);
defparam \top/processor/core_block_363_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_362_s0  (
	.D(\top/processor/block_buffer [362]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [362])
);
defparam \top/processor/core_block_362_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_361_s0  (
	.D(\top/processor/block_buffer [361]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [361])
);
defparam \top/processor/core_block_361_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_360_s0  (
	.D(\top/processor/block_buffer [360]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [360])
);
defparam \top/processor/core_block_360_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_359_s0  (
	.D(\top/processor/block_buffer [359]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [359])
);
defparam \top/processor/core_block_359_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_358_s0  (
	.D(\top/processor/block_buffer [358]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [358])
);
defparam \top/processor/core_block_358_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_357_s0  (
	.D(\top/processor/block_buffer [357]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [357])
);
defparam \top/processor/core_block_357_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_356_s0  (
	.D(\top/processor/block_buffer [356]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [356])
);
defparam \top/processor/core_block_356_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_355_s0  (
	.D(\top/processor/block_buffer [355]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [355])
);
defparam \top/processor/core_block_355_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_354_s0  (
	.D(\top/processor/block_buffer [354]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [354])
);
defparam \top/processor/core_block_354_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_353_s0  (
	.D(\top/processor/block_buffer [353]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [353])
);
defparam \top/processor/core_block_353_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_352_s0  (
	.D(\top/processor/block_buffer [352]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [352])
);
defparam \top/processor/core_block_352_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_351_s0  (
	.D(\top/processor/block_buffer [351]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [351])
);
defparam \top/processor/core_block_351_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_350_s0  (
	.D(\top/processor/block_buffer [350]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [350])
);
defparam \top/processor/core_block_350_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_349_s0  (
	.D(\top/processor/block_buffer [349]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [349])
);
defparam \top/processor/core_block_349_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_348_s0  (
	.D(\top/processor/block_buffer [348]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [348])
);
defparam \top/processor/core_block_348_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_347_s0  (
	.D(\top/processor/block_buffer [347]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [347])
);
defparam \top/processor/core_block_347_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_346_s0  (
	.D(\top/processor/block_buffer [346]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [346])
);
defparam \top/processor/core_block_346_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_345_s0  (
	.D(\top/processor/block_buffer [345]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [345])
);
defparam \top/processor/core_block_345_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_344_s0  (
	.D(\top/processor/block_buffer [344]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [344])
);
defparam \top/processor/core_block_344_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_343_s0  (
	.D(\top/processor/block_buffer [343]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [343])
);
defparam \top/processor/core_block_343_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_342_s0  (
	.D(\top/processor/block_buffer [342]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [342])
);
defparam \top/processor/core_block_342_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_341_s0  (
	.D(\top/processor/block_buffer [341]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [341])
);
defparam \top/processor/core_block_341_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_340_s0  (
	.D(\top/processor/block_buffer [340]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [340])
);
defparam \top/processor/core_block_340_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_339_s0  (
	.D(\top/processor/block_buffer [339]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [339])
);
defparam \top/processor/core_block_339_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_338_s0  (
	.D(\top/processor/block_buffer [338]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [338])
);
defparam \top/processor/core_block_338_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_337_s0  (
	.D(\top/processor/block_buffer [337]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [337])
);
defparam \top/processor/core_block_337_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_336_s0  (
	.D(\top/processor/block_buffer [336]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [336])
);
defparam \top/processor/core_block_336_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_335_s0  (
	.D(\top/processor/block_buffer [335]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [335])
);
defparam \top/processor/core_block_335_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_334_s0  (
	.D(\top/processor/block_buffer [334]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [334])
);
defparam \top/processor/core_block_334_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_333_s0  (
	.D(\top/processor/block_buffer [333]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [333])
);
defparam \top/processor/core_block_333_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_332_s0  (
	.D(\top/processor/block_buffer [332]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [332])
);
defparam \top/processor/core_block_332_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_331_s0  (
	.D(\top/processor/block_buffer [331]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [331])
);
defparam \top/processor/core_block_331_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_330_s0  (
	.D(\top/processor/block_buffer [330]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [330])
);
defparam \top/processor/core_block_330_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_329_s0  (
	.D(\top/processor/block_buffer [329]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [329])
);
defparam \top/processor/core_block_329_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_328_s0  (
	.D(\top/processor/block_buffer [328]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [328])
);
defparam \top/processor/core_block_328_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_327_s0  (
	.D(\top/processor/block_buffer [327]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [327])
);
defparam \top/processor/core_block_327_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_326_s0  (
	.D(\top/processor/block_buffer [326]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [326])
);
defparam \top/processor/core_block_326_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_325_s0  (
	.D(\top/processor/block_buffer [325]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [325])
);
defparam \top/processor/core_block_325_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_324_s0  (
	.D(\top/processor/block_buffer [324]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [324])
);
defparam \top/processor/core_block_324_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_323_s0  (
	.D(\top/processor/block_buffer [323]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [323])
);
defparam \top/processor/core_block_323_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_322_s0  (
	.D(\top/processor/block_buffer [322]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [322])
);
defparam \top/processor/core_block_322_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_321_s0  (
	.D(\top/processor/block_buffer [321]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [321])
);
defparam \top/processor/core_block_321_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_320_s0  (
	.D(\top/processor/block_buffer [320]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [320])
);
defparam \top/processor/core_block_320_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_319_s0  (
	.D(\top/processor/block_buffer [319]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [319])
);
defparam \top/processor/core_block_319_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_318_s0  (
	.D(\top/processor/block_buffer [318]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [318])
);
defparam \top/processor/core_block_318_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_317_s0  (
	.D(\top/processor/block_buffer [317]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [317])
);
defparam \top/processor/core_block_317_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_316_s0  (
	.D(\top/processor/block_buffer [316]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [316])
);
defparam \top/processor/core_block_316_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_315_s0  (
	.D(\top/processor/block_buffer [315]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [315])
);
defparam \top/processor/core_block_315_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_314_s0  (
	.D(\top/processor/block_buffer [314]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [314])
);
defparam \top/processor/core_block_314_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_313_s0  (
	.D(\top/processor/block_buffer [313]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [313])
);
defparam \top/processor/core_block_313_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_312_s0  (
	.D(\top/processor/block_buffer [312]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [312])
);
defparam \top/processor/core_block_312_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_311_s0  (
	.D(\top/processor/block_buffer [311]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [311])
);
defparam \top/processor/core_block_311_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_310_s0  (
	.D(\top/processor/block_buffer [310]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [310])
);
defparam \top/processor/core_block_310_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_309_s0  (
	.D(\top/processor/block_buffer [309]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [309])
);
defparam \top/processor/core_block_309_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_308_s0  (
	.D(\top/processor/block_buffer [308]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [308])
);
defparam \top/processor/core_block_308_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_307_s0  (
	.D(\top/processor/block_buffer [307]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [307])
);
defparam \top/processor/core_block_307_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_306_s0  (
	.D(\top/processor/block_buffer [306]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [306])
);
defparam \top/processor/core_block_306_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_305_s0  (
	.D(\top/processor/block_buffer [305]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [305])
);
defparam \top/processor/core_block_305_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_304_s0  (
	.D(\top/processor/block_buffer [304]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [304])
);
defparam \top/processor/core_block_304_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_303_s0  (
	.D(\top/processor/block_buffer [303]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [303])
);
defparam \top/processor/core_block_303_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_302_s0  (
	.D(\top/processor/block_buffer [302]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [302])
);
defparam \top/processor/core_block_302_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_301_s0  (
	.D(\top/processor/block_buffer [301]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [301])
);
defparam \top/processor/core_block_301_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_300_s0  (
	.D(\top/processor/block_buffer [300]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [300])
);
defparam \top/processor/core_block_300_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_299_s0  (
	.D(\top/processor/block_buffer [299]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [299])
);
defparam \top/processor/core_block_299_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_298_s0  (
	.D(\top/processor/block_buffer [298]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [298])
);
defparam \top/processor/core_block_298_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_297_s0  (
	.D(\top/processor/block_buffer [297]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [297])
);
defparam \top/processor/core_block_297_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_296_s0  (
	.D(\top/processor/block_buffer [296]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [296])
);
defparam \top/processor/core_block_296_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_295_s0  (
	.D(\top/processor/block_buffer [295]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [295])
);
defparam \top/processor/core_block_295_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_294_s0  (
	.D(\top/processor/block_buffer [294]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [294])
);
defparam \top/processor/core_block_294_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_293_s0  (
	.D(\top/processor/block_buffer [293]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [293])
);
defparam \top/processor/core_block_293_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_292_s0  (
	.D(\top/processor/block_buffer [292]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [292])
);
defparam \top/processor/core_block_292_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_291_s0  (
	.D(\top/processor/block_buffer [291]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [291])
);
defparam \top/processor/core_block_291_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_290_s0  (
	.D(\top/processor/block_buffer [290]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [290])
);
defparam \top/processor/core_block_290_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_289_s0  (
	.D(\top/processor/block_buffer [289]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [289])
);
defparam \top/processor/core_block_289_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_288_s0  (
	.D(\top/processor/block_buffer [288]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [288])
);
defparam \top/processor/core_block_288_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_287_s0  (
	.D(\top/processor/block_buffer [287]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [287])
);
defparam \top/processor/core_block_287_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_286_s0  (
	.D(\top/processor/block_buffer [286]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [286])
);
defparam \top/processor/core_block_286_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_285_s0  (
	.D(\top/processor/block_buffer [285]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [285])
);
defparam \top/processor/core_block_285_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_284_s0  (
	.D(\top/processor/block_buffer [284]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [284])
);
defparam \top/processor/core_block_284_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_283_s0  (
	.D(\top/processor/block_buffer [283]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [283])
);
defparam \top/processor/core_block_283_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_282_s0  (
	.D(\top/processor/block_buffer [282]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [282])
);
defparam \top/processor/core_block_282_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_281_s0  (
	.D(\top/processor/block_buffer [281]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [281])
);
defparam \top/processor/core_block_281_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_280_s0  (
	.D(\top/processor/block_buffer [280]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [280])
);
defparam \top/processor/core_block_280_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_279_s0  (
	.D(\top/processor/block_buffer [279]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [279])
);
defparam \top/processor/core_block_279_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_278_s0  (
	.D(\top/processor/block_buffer [278]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [278])
);
defparam \top/processor/core_block_278_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_277_s0  (
	.D(\top/processor/block_buffer [277]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [277])
);
defparam \top/processor/core_block_277_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_276_s0  (
	.D(\top/processor/block_buffer [276]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [276])
);
defparam \top/processor/core_block_276_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_275_s0  (
	.D(\top/processor/block_buffer [275]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [275])
);
defparam \top/processor/core_block_275_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_274_s0  (
	.D(\top/processor/block_buffer [274]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [274])
);
defparam \top/processor/core_block_274_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_273_s0  (
	.D(\top/processor/block_buffer [273]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [273])
);
defparam \top/processor/core_block_273_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_272_s0  (
	.D(\top/processor/block_buffer [272]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [272])
);
defparam \top/processor/core_block_272_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_271_s0  (
	.D(\top/processor/block_buffer [271]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [271])
);
defparam \top/processor/core_block_271_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_270_s0  (
	.D(\top/processor/block_buffer [270]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [270])
);
defparam \top/processor/core_block_270_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_269_s0  (
	.D(\top/processor/block_buffer [269]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [269])
);
defparam \top/processor/core_block_269_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_268_s0  (
	.D(\top/processor/block_buffer [268]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [268])
);
defparam \top/processor/core_block_268_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_267_s0  (
	.D(\top/processor/block_buffer [267]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [267])
);
defparam \top/processor/core_block_267_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_266_s0  (
	.D(\top/processor/block_buffer [266]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [266])
);
defparam \top/processor/core_block_266_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_265_s0  (
	.D(\top/processor/block_buffer [265]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [265])
);
defparam \top/processor/core_block_265_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_264_s0  (
	.D(\top/processor/block_buffer [264]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [264])
);
defparam \top/processor/core_block_264_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_263_s0  (
	.D(\top/processor/block_buffer [263]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [263])
);
defparam \top/processor/core_block_263_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_262_s0  (
	.D(\top/processor/block_buffer [262]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [262])
);
defparam \top/processor/core_block_262_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_261_s0  (
	.D(\top/processor/block_buffer [261]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [261])
);
defparam \top/processor/core_block_261_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_260_s0  (
	.D(\top/processor/block_buffer [260]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [260])
);
defparam \top/processor/core_block_260_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_259_s0  (
	.D(\top/processor/block_buffer [259]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [259])
);
defparam \top/processor/core_block_259_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_258_s0  (
	.D(\top/processor/block_buffer [258]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [258])
);
defparam \top/processor/core_block_258_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_257_s0  (
	.D(\top/processor/block_buffer [257]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [257])
);
defparam \top/processor/core_block_257_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_256_s0  (
	.D(\top/processor/block_buffer [256]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [256])
);
defparam \top/processor/core_block_256_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_255_s0  (
	.D(\top/processor/block_buffer [255]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [255])
);
defparam \top/processor/core_block_255_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_254_s0  (
	.D(\top/processor/block_buffer [254]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [254])
);
defparam \top/processor/core_block_254_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_253_s0  (
	.D(\top/processor/block_buffer [253]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [253])
);
defparam \top/processor/core_block_253_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_252_s0  (
	.D(\top/processor/block_buffer [252]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [252])
);
defparam \top/processor/core_block_252_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_251_s0  (
	.D(\top/processor/block_buffer [251]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [251])
);
defparam \top/processor/core_block_251_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_250_s0  (
	.D(\top/processor/block_buffer [250]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [250])
);
defparam \top/processor/core_block_250_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_249_s0  (
	.D(\top/processor/block_buffer [249]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [249])
);
defparam \top/processor/core_block_249_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_248_s0  (
	.D(\top/processor/block_buffer [248]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [248])
);
defparam \top/processor/core_block_248_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_247_s0  (
	.D(\top/processor/block_buffer [247]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [247])
);
defparam \top/processor/core_block_247_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_246_s0  (
	.D(\top/processor/block_buffer [246]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [246])
);
defparam \top/processor/core_block_246_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_245_s0  (
	.D(\top/processor/block_buffer [245]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [245])
);
defparam \top/processor/core_block_245_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_244_s0  (
	.D(\top/processor/block_buffer [244]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [244])
);
defparam \top/processor/core_block_244_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_243_s0  (
	.D(\top/processor/block_buffer [243]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [243])
);
defparam \top/processor/core_block_243_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_242_s0  (
	.D(\top/processor/block_buffer [242]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [242])
);
defparam \top/processor/core_block_242_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_241_s0  (
	.D(\top/processor/block_buffer [241]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [241])
);
defparam \top/processor/core_block_241_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_240_s0  (
	.D(\top/processor/block_buffer [240]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [240])
);
defparam \top/processor/core_block_240_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_239_s0  (
	.D(\top/processor/block_buffer [239]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [239])
);
defparam \top/processor/core_block_239_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_238_s0  (
	.D(\top/processor/block_buffer [238]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [238])
);
defparam \top/processor/core_block_238_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_237_s0  (
	.D(\top/processor/block_buffer [237]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [237])
);
defparam \top/processor/core_block_237_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_236_s0  (
	.D(\top/processor/block_buffer [236]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [236])
);
defparam \top/processor/core_block_236_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_235_s0  (
	.D(\top/processor/block_buffer [235]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [235])
);
defparam \top/processor/core_block_235_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_234_s0  (
	.D(\top/processor/block_buffer [234]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [234])
);
defparam \top/processor/core_block_234_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_233_s0  (
	.D(\top/processor/block_buffer [233]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [233])
);
defparam \top/processor/core_block_233_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_232_s0  (
	.D(\top/processor/block_buffer [232]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [232])
);
defparam \top/processor/core_block_232_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_231_s0  (
	.D(\top/processor/block_buffer [231]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [231])
);
defparam \top/processor/core_block_231_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_230_s0  (
	.D(\top/processor/block_buffer [230]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [230])
);
defparam \top/processor/core_block_230_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_229_s0  (
	.D(\top/processor/block_buffer [229]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [229])
);
defparam \top/processor/core_block_229_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_228_s0  (
	.D(\top/processor/block_buffer [228]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [228])
);
defparam \top/processor/core_block_228_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_227_s0  (
	.D(\top/processor/block_buffer [227]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [227])
);
defparam \top/processor/core_block_227_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_226_s0  (
	.D(\top/processor/block_buffer [226]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [226])
);
defparam \top/processor/core_block_226_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_225_s0  (
	.D(\top/processor/block_buffer [225]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [225])
);
defparam \top/processor/core_block_225_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_224_s0  (
	.D(\top/processor/block_buffer [224]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [224])
);
defparam \top/processor/core_block_224_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_223_s0  (
	.D(\top/processor/block_buffer [223]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [223])
);
defparam \top/processor/core_block_223_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_222_s0  (
	.D(\top/processor/block_buffer [222]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [222])
);
defparam \top/processor/core_block_222_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_221_s0  (
	.D(\top/processor/block_buffer [221]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [221])
);
defparam \top/processor/core_block_221_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_220_s0  (
	.D(\top/processor/block_buffer [220]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [220])
);
defparam \top/processor/core_block_220_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_219_s0  (
	.D(\top/processor/block_buffer [219]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [219])
);
defparam \top/processor/core_block_219_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_218_s0  (
	.D(\top/processor/block_buffer [218]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [218])
);
defparam \top/processor/core_block_218_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_217_s0  (
	.D(\top/processor/block_buffer [217]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [217])
);
defparam \top/processor/core_block_217_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_216_s0  (
	.D(\top/processor/block_buffer [216]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [216])
);
defparam \top/processor/core_block_216_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_215_s0  (
	.D(\top/processor/block_buffer [215]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [215])
);
defparam \top/processor/core_block_215_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_214_s0  (
	.D(\top/processor/block_buffer [214]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [214])
);
defparam \top/processor/core_block_214_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_213_s0  (
	.D(\top/processor/block_buffer [213]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [213])
);
defparam \top/processor/core_block_213_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_212_s0  (
	.D(\top/processor/block_buffer [212]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [212])
);
defparam \top/processor/core_block_212_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_211_s0  (
	.D(\top/processor/block_buffer [211]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [211])
);
defparam \top/processor/core_block_211_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_210_s0  (
	.D(\top/processor/block_buffer [210]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [210])
);
defparam \top/processor/core_block_210_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_209_s0  (
	.D(\top/processor/block_buffer [209]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [209])
);
defparam \top/processor/core_block_209_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_208_s0  (
	.D(\top/processor/block_buffer [208]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [208])
);
defparam \top/processor/core_block_208_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_207_s0  (
	.D(\top/processor/block_buffer [207]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [207])
);
defparam \top/processor/core_block_207_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_206_s0  (
	.D(\top/processor/block_buffer [206]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [206])
);
defparam \top/processor/core_block_206_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_205_s0  (
	.D(\top/processor/block_buffer [205]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [205])
);
defparam \top/processor/core_block_205_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_204_s0  (
	.D(\top/processor/block_buffer [204]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [204])
);
defparam \top/processor/core_block_204_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_203_s0  (
	.D(\top/processor/block_buffer [203]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [203])
);
defparam \top/processor/core_block_203_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_202_s0  (
	.D(\top/processor/block_buffer [202]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [202])
);
defparam \top/processor/core_block_202_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_201_s0  (
	.D(\top/processor/block_buffer [201]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [201])
);
defparam \top/processor/core_block_201_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_200_s0  (
	.D(\top/processor/block_buffer [200]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [200])
);
defparam \top/processor/core_block_200_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_199_s0  (
	.D(\top/processor/block_buffer [199]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [199])
);
defparam \top/processor/core_block_199_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_198_s0  (
	.D(\top/processor/block_buffer [198]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [198])
);
defparam \top/processor/core_block_198_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_197_s0  (
	.D(\top/processor/block_buffer [197]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [197])
);
defparam \top/processor/core_block_197_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_196_s0  (
	.D(\top/processor/block_buffer [196]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [196])
);
defparam \top/processor/core_block_196_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_195_s0  (
	.D(\top/processor/block_buffer [195]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [195])
);
defparam \top/processor/core_block_195_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_194_s0  (
	.D(\top/processor/block_buffer [194]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [194])
);
defparam \top/processor/core_block_194_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_193_s0  (
	.D(\top/processor/block_buffer [193]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [193])
);
defparam \top/processor/core_block_193_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_192_s0  (
	.D(\top/processor/block_buffer [192]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [192])
);
defparam \top/processor/core_block_192_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_191_s0  (
	.D(\top/processor/block_buffer [191]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [191])
);
defparam \top/processor/core_block_191_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_190_s0  (
	.D(\top/processor/block_buffer [190]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [190])
);
defparam \top/processor/core_block_190_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_189_s0  (
	.D(\top/processor/block_buffer [189]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [189])
);
defparam \top/processor/core_block_189_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_188_s0  (
	.D(\top/processor/block_buffer [188]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [188])
);
defparam \top/processor/core_block_188_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_187_s0  (
	.D(\top/processor/block_buffer [187]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [187])
);
defparam \top/processor/core_block_187_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_186_s0  (
	.D(\top/processor/block_buffer [186]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [186])
);
defparam \top/processor/core_block_186_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_185_s0  (
	.D(\top/processor/block_buffer [185]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [185])
);
defparam \top/processor/core_block_185_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_184_s0  (
	.D(\top/processor/block_buffer [184]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [184])
);
defparam \top/processor/core_block_184_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_183_s0  (
	.D(\top/processor/block_buffer [183]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [183])
);
defparam \top/processor/core_block_183_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_182_s0  (
	.D(\top/processor/block_buffer [182]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [182])
);
defparam \top/processor/core_block_182_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_181_s0  (
	.D(\top/processor/block_buffer [181]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [181])
);
defparam \top/processor/core_block_181_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_180_s0  (
	.D(\top/processor/block_buffer [180]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [180])
);
defparam \top/processor/core_block_180_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_179_s0  (
	.D(\top/processor/block_buffer [179]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [179])
);
defparam \top/processor/core_block_179_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_178_s0  (
	.D(\top/processor/block_buffer [178]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [178])
);
defparam \top/processor/core_block_178_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_177_s0  (
	.D(\top/processor/block_buffer [177]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [177])
);
defparam \top/processor/core_block_177_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_176_s0  (
	.D(\top/processor/block_buffer [176]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [176])
);
defparam \top/processor/core_block_176_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_175_s0  (
	.D(\top/processor/block_buffer [175]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [175])
);
defparam \top/processor/core_block_175_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_174_s0  (
	.D(\top/processor/block_buffer [174]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [174])
);
defparam \top/processor/core_block_174_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_173_s0  (
	.D(\top/processor/block_buffer [173]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [173])
);
defparam \top/processor/core_block_173_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_172_s0  (
	.D(\top/processor/block_buffer [172]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [172])
);
defparam \top/processor/core_block_172_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_171_s0  (
	.D(\top/processor/block_buffer [171]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [171])
);
defparam \top/processor/core_block_171_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_170_s0  (
	.D(\top/processor/block_buffer [170]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [170])
);
defparam \top/processor/core_block_170_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_169_s0  (
	.D(\top/processor/block_buffer [169]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [169])
);
defparam \top/processor/core_block_169_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_168_s0  (
	.D(\top/processor/block_buffer [168]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [168])
);
defparam \top/processor/core_block_168_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_167_s0  (
	.D(\top/processor/block_buffer [167]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [167])
);
defparam \top/processor/core_block_167_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_166_s0  (
	.D(\top/processor/block_buffer [166]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [166])
);
defparam \top/processor/core_block_166_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_165_s0  (
	.D(\top/processor/block_buffer [165]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [165])
);
defparam \top/processor/core_block_165_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_164_s0  (
	.D(\top/processor/block_buffer [164]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [164])
);
defparam \top/processor/core_block_164_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_163_s0  (
	.D(\top/processor/block_buffer [163]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [163])
);
defparam \top/processor/core_block_163_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_162_s0  (
	.D(\top/processor/block_buffer [162]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [162])
);
defparam \top/processor/core_block_162_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_161_s0  (
	.D(\top/processor/block_buffer [161]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [161])
);
defparam \top/processor/core_block_161_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_160_s0  (
	.D(\top/processor/block_buffer [160]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [160])
);
defparam \top/processor/core_block_160_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_159_s0  (
	.D(\top/processor/block_buffer [159]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [159])
);
defparam \top/processor/core_block_159_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_158_s0  (
	.D(\top/processor/block_buffer [158]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [158])
);
defparam \top/processor/core_block_158_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_157_s0  (
	.D(\top/processor/block_buffer [157]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [157])
);
defparam \top/processor/core_block_157_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_156_s0  (
	.D(\top/processor/block_buffer [156]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [156])
);
defparam \top/processor/core_block_156_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_155_s0  (
	.D(\top/processor/block_buffer [155]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [155])
);
defparam \top/processor/core_block_155_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_154_s0  (
	.D(\top/processor/block_buffer [154]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [154])
);
defparam \top/processor/core_block_154_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_153_s0  (
	.D(\top/processor/block_buffer [153]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [153])
);
defparam \top/processor/core_block_153_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_152_s0  (
	.D(\top/processor/block_buffer [152]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [152])
);
defparam \top/processor/core_block_152_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_151_s0  (
	.D(\top/processor/block_buffer [151]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [151])
);
defparam \top/processor/core_block_151_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_150_s0  (
	.D(\top/processor/block_buffer [150]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [150])
);
defparam \top/processor/core_block_150_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_149_s0  (
	.D(\top/processor/block_buffer [149]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [149])
);
defparam \top/processor/core_block_149_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_148_s0  (
	.D(\top/processor/block_buffer [148]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [148])
);
defparam \top/processor/core_block_148_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_147_s0  (
	.D(\top/processor/block_buffer [147]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [147])
);
defparam \top/processor/core_block_147_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_146_s0  (
	.D(\top/processor/block_buffer [146]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [146])
);
defparam \top/processor/core_block_146_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_145_s0  (
	.D(\top/processor/block_buffer [145]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [145])
);
defparam \top/processor/core_block_145_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_144_s0  (
	.D(\top/processor/block_buffer [144]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [144])
);
defparam \top/processor/core_block_144_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_143_s0  (
	.D(\top/processor/block_buffer [143]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [143])
);
defparam \top/processor/core_block_143_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_142_s0  (
	.D(\top/processor/block_buffer [142]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [142])
);
defparam \top/processor/core_block_142_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_141_s0  (
	.D(\top/processor/block_buffer [141]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [141])
);
defparam \top/processor/core_block_141_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_140_s0  (
	.D(\top/processor/block_buffer [140]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [140])
);
defparam \top/processor/core_block_140_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_139_s0  (
	.D(\top/processor/block_buffer [139]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [139])
);
defparam \top/processor/core_block_139_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_138_s0  (
	.D(\top/processor/block_buffer [138]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [138])
);
defparam \top/processor/core_block_138_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_137_s0  (
	.D(\top/processor/block_buffer [137]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [137])
);
defparam \top/processor/core_block_137_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_136_s0  (
	.D(\top/processor/block_buffer [136]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [136])
);
defparam \top/processor/core_block_136_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_135_s0  (
	.D(\top/processor/block_buffer [135]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [135])
);
defparam \top/processor/core_block_135_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_134_s0  (
	.D(\top/processor/block_buffer [134]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [134])
);
defparam \top/processor/core_block_134_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_133_s0  (
	.D(\top/processor/block_buffer [133]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [133])
);
defparam \top/processor/core_block_133_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_132_s0  (
	.D(\top/processor/block_buffer [132]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [132])
);
defparam \top/processor/core_block_132_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_131_s0  (
	.D(\top/processor/block_buffer [131]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [131])
);
defparam \top/processor/core_block_131_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_130_s0  (
	.D(\top/processor/block_buffer [130]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [130])
);
defparam \top/processor/core_block_130_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_129_s0  (
	.D(\top/processor/block_buffer [129]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [129])
);
defparam \top/processor/core_block_129_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_128_s0  (
	.D(\top/processor/block_buffer [128]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [128])
);
defparam \top/processor/core_block_128_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_127_s0  (
	.D(\top/processor/block_buffer [127]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [127])
);
defparam \top/processor/core_block_127_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_126_s0  (
	.D(\top/processor/block_buffer [126]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [126])
);
defparam \top/processor/core_block_126_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_125_s0  (
	.D(\top/processor/block_buffer [125]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [125])
);
defparam \top/processor/core_block_125_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_124_s0  (
	.D(\top/processor/block_buffer [124]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [124])
);
defparam \top/processor/core_block_124_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_123_s0  (
	.D(\top/processor/block_buffer [123]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [123])
);
defparam \top/processor/core_block_123_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_122_s0  (
	.D(\top/processor/block_buffer [122]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [122])
);
defparam \top/processor/core_block_122_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_121_s0  (
	.D(\top/processor/block_buffer [121]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [121])
);
defparam \top/processor/core_block_121_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_120_s0  (
	.D(\top/processor/block_buffer [120]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [120])
);
defparam \top/processor/core_block_120_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_119_s0  (
	.D(\top/processor/block_buffer [119]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [119])
);
defparam \top/processor/core_block_119_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_118_s0  (
	.D(\top/processor/block_buffer [118]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [118])
);
defparam \top/processor/core_block_118_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_117_s0  (
	.D(\top/processor/block_buffer [117]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [117])
);
defparam \top/processor/core_block_117_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_116_s0  (
	.D(\top/processor/block_buffer [116]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [116])
);
defparam \top/processor/core_block_116_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_115_s0  (
	.D(\top/processor/block_buffer [115]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [115])
);
defparam \top/processor/core_block_115_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_114_s0  (
	.D(\top/processor/block_buffer [114]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [114])
);
defparam \top/processor/core_block_114_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_113_s0  (
	.D(\top/processor/block_buffer [113]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [113])
);
defparam \top/processor/core_block_113_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_112_s0  (
	.D(\top/processor/block_buffer [112]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [112])
);
defparam \top/processor/core_block_112_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_111_s0  (
	.D(\top/processor/block_buffer [111]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [111])
);
defparam \top/processor/core_block_111_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_110_s0  (
	.D(\top/processor/block_buffer [110]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [110])
);
defparam \top/processor/core_block_110_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_109_s0  (
	.D(\top/processor/block_buffer [109]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [109])
);
defparam \top/processor/core_block_109_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_108_s0  (
	.D(\top/processor/block_buffer [108]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [108])
);
defparam \top/processor/core_block_108_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_107_s0  (
	.D(\top/processor/block_buffer [107]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [107])
);
defparam \top/processor/core_block_107_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_106_s0  (
	.D(\top/processor/block_buffer [106]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [106])
);
defparam \top/processor/core_block_106_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_105_s0  (
	.D(\top/processor/block_buffer [105]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [105])
);
defparam \top/processor/core_block_105_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_104_s0  (
	.D(\top/processor/block_buffer [104]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [104])
);
defparam \top/processor/core_block_104_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_103_s0  (
	.D(\top/processor/block_buffer [103]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [103])
);
defparam \top/processor/core_block_103_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_102_s0  (
	.D(\top/processor/block_buffer [102]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [102])
);
defparam \top/processor/core_block_102_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_101_s0  (
	.D(\top/processor/block_buffer [101]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [101])
);
defparam \top/processor/core_block_101_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_100_s0  (
	.D(\top/processor/block_buffer [100]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [100])
);
defparam \top/processor/core_block_100_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_99_s0  (
	.D(\top/processor/block_buffer [99]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [99])
);
defparam \top/processor/core_block_99_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_98_s0  (
	.D(\top/processor/block_buffer [98]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [98])
);
defparam \top/processor/core_block_98_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_97_s0  (
	.D(\top/processor/block_buffer [97]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [97])
);
defparam \top/processor/core_block_97_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_96_s0  (
	.D(\top/processor/block_buffer [96]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [96])
);
defparam \top/processor/core_block_96_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_95_s0  (
	.D(\top/processor/block_buffer [95]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [95])
);
defparam \top/processor/core_block_95_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_94_s0  (
	.D(\top/processor/block_buffer [94]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [94])
);
defparam \top/processor/core_block_94_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_93_s0  (
	.D(\top/processor/block_buffer [93]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [93])
);
defparam \top/processor/core_block_93_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_92_s0  (
	.D(\top/processor/block_buffer [92]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [92])
);
defparam \top/processor/core_block_92_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_91_s0  (
	.D(\top/processor/block_buffer [91]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [91])
);
defparam \top/processor/core_block_91_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_90_s0  (
	.D(\top/processor/block_buffer [90]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [90])
);
defparam \top/processor/core_block_90_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_89_s0  (
	.D(\top/processor/block_buffer [89]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [89])
);
defparam \top/processor/core_block_89_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_88_s0  (
	.D(\top/processor/block_buffer [88]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [88])
);
defparam \top/processor/core_block_88_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_87_s0  (
	.D(\top/processor/block_buffer [87]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [87])
);
defparam \top/processor/core_block_87_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_86_s0  (
	.D(\top/processor/block_buffer [86]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [86])
);
defparam \top/processor/core_block_86_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_85_s0  (
	.D(\top/processor/block_buffer [85]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [85])
);
defparam \top/processor/core_block_85_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_84_s0  (
	.D(\top/processor/block_buffer [84]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [84])
);
defparam \top/processor/core_block_84_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_83_s0  (
	.D(\top/processor/block_buffer [83]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [83])
);
defparam \top/processor/core_block_83_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_82_s0  (
	.D(\top/processor/block_buffer [82]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [82])
);
defparam \top/processor/core_block_82_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_81_s0  (
	.D(\top/processor/block_buffer [81]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [81])
);
defparam \top/processor/core_block_81_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_80_s0  (
	.D(\top/processor/block_buffer [80]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [80])
);
defparam \top/processor/core_block_80_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_79_s0  (
	.D(\top/processor/block_buffer [79]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [79])
);
defparam \top/processor/core_block_79_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_78_s0  (
	.D(\top/processor/block_buffer [78]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [78])
);
defparam \top/processor/core_block_78_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_77_s0  (
	.D(\top/processor/block_buffer [77]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [77])
);
defparam \top/processor/core_block_77_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_76_s0  (
	.D(\top/processor/block_buffer [76]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [76])
);
defparam \top/processor/core_block_76_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_75_s0  (
	.D(\top/processor/block_buffer [75]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [75])
);
defparam \top/processor/core_block_75_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_74_s0  (
	.D(\top/processor/block_buffer [74]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [74])
);
defparam \top/processor/core_block_74_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_73_s0  (
	.D(\top/processor/block_buffer [73]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [73])
);
defparam \top/processor/core_block_73_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_72_s0  (
	.D(\top/processor/block_buffer [72]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [72])
);
defparam \top/processor/core_block_72_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_71_s0  (
	.D(\top/processor/block_buffer [71]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [71])
);
defparam \top/processor/core_block_71_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_70_s0  (
	.D(\top/processor/block_buffer [70]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [70])
);
defparam \top/processor/core_block_70_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_69_s0  (
	.D(\top/processor/block_buffer [69]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [69])
);
defparam \top/processor/core_block_69_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_68_s0  (
	.D(\top/processor/block_buffer [68]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [68])
);
defparam \top/processor/core_block_68_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_67_s0  (
	.D(\top/processor/block_buffer [67]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [67])
);
defparam \top/processor/core_block_67_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_66_s0  (
	.D(\top/processor/block_buffer [66]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [66])
);
defparam \top/processor/core_block_66_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_65_s0  (
	.D(\top/processor/block_buffer [65]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [65])
);
defparam \top/processor/core_block_65_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_64_s0  (
	.D(\top/processor/block_buffer [64]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [64])
);
defparam \top/processor/core_block_64_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_63_s0  (
	.D(\top/processor/block_buffer [63]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [63])
);
defparam \top/processor/core_block_63_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_62_s0  (
	.D(\top/processor/block_buffer [62]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [62])
);
defparam \top/processor/core_block_62_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_61_s0  (
	.D(\top/processor/block_buffer [61]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [61])
);
defparam \top/processor/core_block_61_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_60_s0  (
	.D(\top/processor/block_buffer [60]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [60])
);
defparam \top/processor/core_block_60_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_59_s0  (
	.D(\top/processor/block_buffer [59]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [59])
);
defparam \top/processor/core_block_59_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_58_s0  (
	.D(\top/processor/block_buffer [58]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [58])
);
defparam \top/processor/core_block_58_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_57_s0  (
	.D(\top/processor/block_buffer [57]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [57])
);
defparam \top/processor/core_block_57_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_56_s0  (
	.D(\top/processor/block_buffer [56]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [56])
);
defparam \top/processor/core_block_56_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_55_s0  (
	.D(\top/processor/block_buffer [55]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [55])
);
defparam \top/processor/core_block_55_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_54_s0  (
	.D(\top/processor/block_buffer [54]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [54])
);
defparam \top/processor/core_block_54_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_53_s0  (
	.D(\top/processor/block_buffer [53]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [53])
);
defparam \top/processor/core_block_53_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_52_s0  (
	.D(\top/processor/block_buffer [52]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [52])
);
defparam \top/processor/core_block_52_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_51_s0  (
	.D(\top/processor/block_buffer [51]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [51])
);
defparam \top/processor/core_block_51_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_50_s0  (
	.D(\top/processor/block_buffer [50]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [50])
);
defparam \top/processor/core_block_50_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_49_s0  (
	.D(\top/processor/block_buffer [49]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [49])
);
defparam \top/processor/core_block_49_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_48_s0  (
	.D(\top/processor/block_buffer [48]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [48])
);
defparam \top/processor/core_block_48_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_47_s0  (
	.D(\top/processor/block_buffer [47]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [47])
);
defparam \top/processor/core_block_47_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_46_s0  (
	.D(\top/processor/block_buffer [46]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [46])
);
defparam \top/processor/core_block_46_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_45_s0  (
	.D(\top/processor/block_buffer [45]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [45])
);
defparam \top/processor/core_block_45_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_44_s0  (
	.D(\top/processor/block_buffer [44]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [44])
);
defparam \top/processor/core_block_44_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_43_s0  (
	.D(\top/processor/block_buffer [43]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [43])
);
defparam \top/processor/core_block_43_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_42_s0  (
	.D(\top/processor/block_buffer [42]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [42])
);
defparam \top/processor/core_block_42_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_41_s0  (
	.D(\top/processor/block_buffer [41]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [41])
);
defparam \top/processor/core_block_41_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_40_s0  (
	.D(\top/processor/block_buffer [40]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [40])
);
defparam \top/processor/core_block_40_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_39_s0  (
	.D(\top/processor/block_buffer [39]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [39])
);
defparam \top/processor/core_block_39_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_38_s0  (
	.D(\top/processor/block_buffer [38]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [38])
);
defparam \top/processor/core_block_38_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_37_s0  (
	.D(\top/processor/block_buffer [37]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [37])
);
defparam \top/processor/core_block_37_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_36_s0  (
	.D(\top/processor/block_buffer [36]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [36])
);
defparam \top/processor/core_block_36_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_35_s0  (
	.D(\top/processor/block_buffer [35]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [35])
);
defparam \top/processor/core_block_35_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_34_s0  (
	.D(\top/processor/block_buffer [34]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [34])
);
defparam \top/processor/core_block_34_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_33_s0  (
	.D(\top/processor/block_buffer [33]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [33])
);
defparam \top/processor/core_block_33_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_32_s0  (
	.D(\top/processor/block_buffer [32]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [32])
);
defparam \top/processor/core_block_32_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_31_s0  (
	.D(\top/processor/block_buffer [31]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [31])
);
defparam \top/processor/core_block_31_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_30_s0  (
	.D(\top/processor/block_buffer [30]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [30])
);
defparam \top/processor/core_block_30_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_29_s0  (
	.D(\top/processor/block_buffer [29]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [29])
);
defparam \top/processor/core_block_29_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_28_s0  (
	.D(\top/processor/block_buffer [28]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [28])
);
defparam \top/processor/core_block_28_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_27_s0  (
	.D(\top/processor/block_buffer [27]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [27])
);
defparam \top/processor/core_block_27_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_26_s0  (
	.D(\top/processor/block_buffer [26]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [26])
);
defparam \top/processor/core_block_26_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_25_s0  (
	.D(\top/processor/block_buffer [25]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [25])
);
defparam \top/processor/core_block_25_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_24_s0  (
	.D(\top/processor/block_buffer [24]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [24])
);
defparam \top/processor/core_block_24_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_23_s0  (
	.D(\top/processor/block_buffer [23]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [23])
);
defparam \top/processor/core_block_23_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_22_s0  (
	.D(\top/processor/block_buffer [22]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [22])
);
defparam \top/processor/core_block_22_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_21_s0  (
	.D(\top/processor/block_buffer [21]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [21])
);
defparam \top/processor/core_block_21_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_20_s0  (
	.D(\top/processor/block_buffer [20]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [20])
);
defparam \top/processor/core_block_20_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_19_s0  (
	.D(\top/processor/block_buffer [19]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [19])
);
defparam \top/processor/core_block_19_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_18_s0  (
	.D(\top/processor/block_buffer [18]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [18])
);
defparam \top/processor/core_block_18_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_17_s0  (
	.D(\top/processor/block_buffer [17]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [17])
);
defparam \top/processor/core_block_17_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_16_s0  (
	.D(\top/processor/block_buffer [16]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [16])
);
defparam \top/processor/core_block_16_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_15_s0  (
	.D(\top/processor/block_buffer [15]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [15])
);
defparam \top/processor/core_block_15_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_14_s0  (
	.D(\top/processor/block_buffer [14]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [14])
);
defparam \top/processor/core_block_14_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_13_s0  (
	.D(\top/processor/block_buffer [13]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [13])
);
defparam \top/processor/core_block_13_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_12_s0  (
	.D(\top/processor/block_buffer [12]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [12])
);
defparam \top/processor/core_block_12_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_11_s0  (
	.D(\top/processor/block_buffer [11]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [11])
);
defparam \top/processor/core_block_11_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_10_s0  (
	.D(\top/processor/block_buffer [10]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [10])
);
defparam \top/processor/core_block_10_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_9_s0  (
	.D(\top/processor/block_buffer [9]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [9])
);
defparam \top/processor/core_block_9_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_8_s0  (
	.D(\top/processor/block_buffer [8]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [8])
);
defparam \top/processor/core_block_8_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_7_s0  (
	.D(\top/processor/block_buffer [7]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [7])
);
defparam \top/processor/core_block_7_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_6_s0  (
	.D(\top/processor/block_buffer [6]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [6])
);
defparam \top/processor/core_block_6_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_5_s0  (
	.D(\top/processor/block_buffer [5]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [5])
);
defparam \top/processor/core_block_5_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_4_s0  (
	.D(\top/processor/block_buffer [4]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [4])
);
defparam \top/processor/core_block_4_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_3_s0  (
	.D(\top/processor/block_buffer [3]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [3])
);
defparam \top/processor/core_block_3_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_2_s0  (
	.D(\top/processor/block_buffer [2]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [2])
);
defparam \top/processor/core_block_2_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_1_s0  (
	.D(\top/processor/block_buffer [1]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [1])
);
defparam \top/processor/core_block_1_s0 .INIT=1'b0;
DFFCE \top/processor/core_block_0_s0  (
	.D(\top/processor/block_buffer [0]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_block [0])
);
defparam \top/processor/core_block_0_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_255_s0  (
	.D(\top/hash_out [255]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [255])
);
defparam \top/processor/core_hash_init_255_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_254_s0  (
	.D(\top/hash_out [254]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [254])
);
defparam \top/processor/core_hash_init_254_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_253_s0  (
	.D(\top/hash_out [253]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [253])
);
defparam \top/processor/core_hash_init_253_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_252_s0  (
	.D(\top/hash_out [252]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [252])
);
defparam \top/processor/core_hash_init_252_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_251_s0  (
	.D(\top/hash_out [251]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [251])
);
defparam \top/processor/core_hash_init_251_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_250_s0  (
	.D(\top/hash_out [250]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [250])
);
defparam \top/processor/core_hash_init_250_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_249_s0  (
	.D(\top/hash_out [249]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [249])
);
defparam \top/processor/core_hash_init_249_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_248_s0  (
	.D(\top/hash_out [248]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [248])
);
defparam \top/processor/core_hash_init_248_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_247_s0  (
	.D(\top/hash_out [247]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [247])
);
defparam \top/processor/core_hash_init_247_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_246_s0  (
	.D(\top/hash_out [246]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [246])
);
defparam \top/processor/core_hash_init_246_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_245_s0  (
	.D(\top/hash_out [245]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [245])
);
defparam \top/processor/core_hash_init_245_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_244_s0  (
	.D(\top/hash_out [244]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [244])
);
defparam \top/processor/core_hash_init_244_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_243_s0  (
	.D(\top/hash_out [243]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [243])
);
defparam \top/processor/core_hash_init_243_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_242_s0  (
	.D(\top/hash_out [242]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [242])
);
defparam \top/processor/core_hash_init_242_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_241_s0  (
	.D(\top/hash_out [241]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [241])
);
defparam \top/processor/core_hash_init_241_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_240_s0  (
	.D(\top/hash_out [240]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [240])
);
defparam \top/processor/core_hash_init_240_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_239_s0  (
	.D(\top/hash_out [239]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [239])
);
defparam \top/processor/core_hash_init_239_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_238_s0  (
	.D(\top/hash_out [238]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [238])
);
defparam \top/processor/core_hash_init_238_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_237_s0  (
	.D(\top/hash_out [237]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [237])
);
defparam \top/processor/core_hash_init_237_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_236_s0  (
	.D(\top/hash_out [236]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [236])
);
defparam \top/processor/core_hash_init_236_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_235_s0  (
	.D(\top/hash_out [235]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [235])
);
defparam \top/processor/core_hash_init_235_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_234_s0  (
	.D(\top/hash_out [234]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [234])
);
defparam \top/processor/core_hash_init_234_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_233_s0  (
	.D(\top/hash_out [233]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [233])
);
defparam \top/processor/core_hash_init_233_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_232_s0  (
	.D(\top/hash_out [232]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [232])
);
defparam \top/processor/core_hash_init_232_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_231_s0  (
	.D(\top/hash_out [231]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [231])
);
defparam \top/processor/core_hash_init_231_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_230_s0  (
	.D(\top/hash_out [230]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [230])
);
defparam \top/processor/core_hash_init_230_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_229_s0  (
	.D(\top/hash_out [229]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [229])
);
defparam \top/processor/core_hash_init_229_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_228_s0  (
	.D(\top/hash_out [228]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [228])
);
defparam \top/processor/core_hash_init_228_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_227_s0  (
	.D(\top/hash_out [227]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [227])
);
defparam \top/processor/core_hash_init_227_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_226_s0  (
	.D(\top/hash_out [226]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [226])
);
defparam \top/processor/core_hash_init_226_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_225_s0  (
	.D(\top/hash_out [225]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [225])
);
defparam \top/processor/core_hash_init_225_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_224_s0  (
	.D(\top/hash_out [224]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [224])
);
defparam \top/processor/core_hash_init_224_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_223_s0  (
	.D(\top/hash_out [223]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [223])
);
defparam \top/processor/core_hash_init_223_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_222_s0  (
	.D(\top/hash_out [222]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [222])
);
defparam \top/processor/core_hash_init_222_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_221_s0  (
	.D(\top/hash_out [221]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [221])
);
defparam \top/processor/core_hash_init_221_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_220_s0  (
	.D(\top/hash_out [220]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [220])
);
defparam \top/processor/core_hash_init_220_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_219_s0  (
	.D(\top/hash_out [219]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [219])
);
defparam \top/processor/core_hash_init_219_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_218_s0  (
	.D(\top/hash_out [218]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [218])
);
defparam \top/processor/core_hash_init_218_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_217_s0  (
	.D(\top/hash_out [217]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [217])
);
defparam \top/processor/core_hash_init_217_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_216_s0  (
	.D(\top/hash_out [216]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [216])
);
defparam \top/processor/core_hash_init_216_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_215_s0  (
	.D(\top/hash_out [215]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [215])
);
defparam \top/processor/core_hash_init_215_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_214_s0  (
	.D(\top/hash_out [214]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [214])
);
defparam \top/processor/core_hash_init_214_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_213_s0  (
	.D(\top/hash_out [213]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [213])
);
defparam \top/processor/core_hash_init_213_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_212_s0  (
	.D(\top/hash_out [212]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [212])
);
defparam \top/processor/core_hash_init_212_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_211_s0  (
	.D(\top/hash_out [211]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [211])
);
defparam \top/processor/core_hash_init_211_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_210_s0  (
	.D(\top/hash_out [210]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [210])
);
defparam \top/processor/core_hash_init_210_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_209_s0  (
	.D(\top/hash_out [209]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [209])
);
defparam \top/processor/core_hash_init_209_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_208_s0  (
	.D(\top/hash_out [208]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [208])
);
defparam \top/processor/core_hash_init_208_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_207_s0  (
	.D(\top/hash_out [207]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [207])
);
defparam \top/processor/core_hash_init_207_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_206_s0  (
	.D(\top/hash_out [206]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [206])
);
defparam \top/processor/core_hash_init_206_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_205_s0  (
	.D(\top/hash_out [205]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [205])
);
defparam \top/processor/core_hash_init_205_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_204_s0  (
	.D(\top/hash_out [204]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [204])
);
defparam \top/processor/core_hash_init_204_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_203_s0  (
	.D(\top/hash_out [203]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [203])
);
defparam \top/processor/core_hash_init_203_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_202_s0  (
	.D(\top/hash_out [202]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [202])
);
defparam \top/processor/core_hash_init_202_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_201_s0  (
	.D(\top/hash_out [201]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [201])
);
defparam \top/processor/core_hash_init_201_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_200_s0  (
	.D(\top/hash_out [200]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [200])
);
defparam \top/processor/core_hash_init_200_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_199_s0  (
	.D(\top/hash_out [199]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [199])
);
defparam \top/processor/core_hash_init_199_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_198_s0  (
	.D(\top/hash_out [198]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [198])
);
defparam \top/processor/core_hash_init_198_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_197_s0  (
	.D(\top/hash_out [197]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [197])
);
defparam \top/processor/core_hash_init_197_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_196_s0  (
	.D(\top/hash_out [196]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [196])
);
defparam \top/processor/core_hash_init_196_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_195_s0  (
	.D(\top/hash_out [195]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [195])
);
defparam \top/processor/core_hash_init_195_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_194_s0  (
	.D(\top/hash_out [194]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [194])
);
defparam \top/processor/core_hash_init_194_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_193_s0  (
	.D(\top/hash_out [193]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [193])
);
defparam \top/processor/core_hash_init_193_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_192_s0  (
	.D(\top/hash_out [192]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [192])
);
defparam \top/processor/core_hash_init_192_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_191_s0  (
	.D(\top/hash_out [191]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [191])
);
defparam \top/processor/core_hash_init_191_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_190_s0  (
	.D(\top/hash_out [190]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [190])
);
defparam \top/processor/core_hash_init_190_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_189_s0  (
	.D(\top/hash_out [189]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [189])
);
defparam \top/processor/core_hash_init_189_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_188_s0  (
	.D(\top/hash_out [188]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [188])
);
defparam \top/processor/core_hash_init_188_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_187_s0  (
	.D(\top/hash_out [187]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [187])
);
defparam \top/processor/core_hash_init_187_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_186_s0  (
	.D(\top/hash_out [186]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [186])
);
defparam \top/processor/core_hash_init_186_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_185_s0  (
	.D(\top/hash_out [185]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [185])
);
defparam \top/processor/core_hash_init_185_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_184_s0  (
	.D(\top/hash_out [184]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [184])
);
defparam \top/processor/core_hash_init_184_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_183_s0  (
	.D(\top/hash_out [183]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [183])
);
defparam \top/processor/core_hash_init_183_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_182_s0  (
	.D(\top/hash_out [182]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [182])
);
defparam \top/processor/core_hash_init_182_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_181_s0  (
	.D(\top/hash_out [181]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [181])
);
defparam \top/processor/core_hash_init_181_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_180_s0  (
	.D(\top/hash_out [180]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [180])
);
defparam \top/processor/core_hash_init_180_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_179_s0  (
	.D(\top/hash_out [179]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [179])
);
defparam \top/processor/core_hash_init_179_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_178_s0  (
	.D(\top/hash_out [178]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [178])
);
defparam \top/processor/core_hash_init_178_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_177_s0  (
	.D(\top/hash_out [177]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [177])
);
defparam \top/processor/core_hash_init_177_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_176_s0  (
	.D(\top/hash_out [176]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [176])
);
defparam \top/processor/core_hash_init_176_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_175_s0  (
	.D(\top/hash_out [175]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [175])
);
defparam \top/processor/core_hash_init_175_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_174_s0  (
	.D(\top/hash_out [174]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [174])
);
defparam \top/processor/core_hash_init_174_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_173_s0  (
	.D(\top/hash_out [173]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [173])
);
defparam \top/processor/core_hash_init_173_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_172_s0  (
	.D(\top/hash_out [172]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [172])
);
defparam \top/processor/core_hash_init_172_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_171_s0  (
	.D(\top/hash_out [171]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [171])
);
defparam \top/processor/core_hash_init_171_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_170_s0  (
	.D(\top/hash_out [170]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [170])
);
defparam \top/processor/core_hash_init_170_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_169_s0  (
	.D(\top/hash_out [169]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [169])
);
defparam \top/processor/core_hash_init_169_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_168_s0  (
	.D(\top/hash_out [168]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [168])
);
defparam \top/processor/core_hash_init_168_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_167_s0  (
	.D(\top/hash_out [167]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [167])
);
defparam \top/processor/core_hash_init_167_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_166_s0  (
	.D(\top/hash_out [166]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [166])
);
defparam \top/processor/core_hash_init_166_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_165_s0  (
	.D(\top/hash_out [165]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [165])
);
defparam \top/processor/core_hash_init_165_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_164_s0  (
	.D(\top/hash_out [164]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [164])
);
defparam \top/processor/core_hash_init_164_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_163_s0  (
	.D(\top/hash_out [163]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [163])
);
defparam \top/processor/core_hash_init_163_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_162_s0  (
	.D(\top/hash_out [162]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [162])
);
defparam \top/processor/core_hash_init_162_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_161_s0  (
	.D(\top/hash_out [161]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [161])
);
defparam \top/processor/core_hash_init_161_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_160_s0  (
	.D(\top/hash_out [160]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [160])
);
defparam \top/processor/core_hash_init_160_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_159_s0  (
	.D(\top/hash_out [159]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [159])
);
defparam \top/processor/core_hash_init_159_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_158_s0  (
	.D(\top/hash_out [158]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [158])
);
defparam \top/processor/core_hash_init_158_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_157_s0  (
	.D(\top/hash_out [157]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [157])
);
defparam \top/processor/core_hash_init_157_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_156_s0  (
	.D(\top/hash_out [156]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [156])
);
defparam \top/processor/core_hash_init_156_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_155_s0  (
	.D(\top/hash_out [155]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [155])
);
defparam \top/processor/core_hash_init_155_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_154_s0  (
	.D(\top/hash_out [154]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [154])
);
defparam \top/processor/core_hash_init_154_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_153_s0  (
	.D(\top/hash_out [153]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [153])
);
defparam \top/processor/core_hash_init_153_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_152_s0  (
	.D(\top/hash_out [152]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [152])
);
defparam \top/processor/core_hash_init_152_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_151_s0  (
	.D(\top/hash_out [151]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [151])
);
defparam \top/processor/core_hash_init_151_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_150_s0  (
	.D(\top/hash_out [150]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [150])
);
defparam \top/processor/core_hash_init_150_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_149_s0  (
	.D(\top/hash_out [149]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [149])
);
defparam \top/processor/core_hash_init_149_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_148_s0  (
	.D(\top/hash_out [148]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [148])
);
defparam \top/processor/core_hash_init_148_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_147_s0  (
	.D(\top/hash_out [147]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [147])
);
defparam \top/processor/core_hash_init_147_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_146_s0  (
	.D(\top/hash_out [146]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [146])
);
defparam \top/processor/core_hash_init_146_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_145_s0  (
	.D(\top/hash_out [145]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [145])
);
defparam \top/processor/core_hash_init_145_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_144_s0  (
	.D(\top/hash_out [144]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [144])
);
defparam \top/processor/core_hash_init_144_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_143_s0  (
	.D(\top/hash_out [143]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [143])
);
defparam \top/processor/core_hash_init_143_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_142_s0  (
	.D(\top/hash_out [142]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [142])
);
defparam \top/processor/core_hash_init_142_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_141_s0  (
	.D(\top/hash_out [141]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [141])
);
defparam \top/processor/core_hash_init_141_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_140_s0  (
	.D(\top/hash_out [140]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [140])
);
defparam \top/processor/core_hash_init_140_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_139_s0  (
	.D(\top/hash_out [139]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [139])
);
defparam \top/processor/core_hash_init_139_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_138_s0  (
	.D(\top/hash_out [138]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [138])
);
defparam \top/processor/core_hash_init_138_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_137_s0  (
	.D(\top/hash_out [137]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [137])
);
defparam \top/processor/core_hash_init_137_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_136_s0  (
	.D(\top/hash_out [136]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [136])
);
defparam \top/processor/core_hash_init_136_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_135_s0  (
	.D(\top/hash_out [135]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [135])
);
defparam \top/processor/core_hash_init_135_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_134_s0  (
	.D(\top/hash_out [134]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [134])
);
defparam \top/processor/core_hash_init_134_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_133_s0  (
	.D(\top/hash_out [133]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [133])
);
defparam \top/processor/core_hash_init_133_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_132_s0  (
	.D(\top/hash_out [132]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [132])
);
defparam \top/processor/core_hash_init_132_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_131_s0  (
	.D(\top/hash_out [131]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [131])
);
defparam \top/processor/core_hash_init_131_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_130_s0  (
	.D(\top/hash_out [130]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [130])
);
defparam \top/processor/core_hash_init_130_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_129_s0  (
	.D(\top/hash_out [129]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [129])
);
defparam \top/processor/core_hash_init_129_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_128_s0  (
	.D(\top/hash_out [128]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [128])
);
defparam \top/processor/core_hash_init_128_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_127_s0  (
	.D(\top/hash_out [127]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [127])
);
defparam \top/processor/core_hash_init_127_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_126_s0  (
	.D(\top/hash_out [126]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [126])
);
defparam \top/processor/core_hash_init_126_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_125_s0  (
	.D(\top/hash_out [125]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [125])
);
defparam \top/processor/core_hash_init_125_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_124_s0  (
	.D(\top/hash_out [124]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [124])
);
defparam \top/processor/core_hash_init_124_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_123_s0  (
	.D(\top/hash_out [123]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [123])
);
defparam \top/processor/core_hash_init_123_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_122_s0  (
	.D(\top/hash_out [122]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [122])
);
defparam \top/processor/core_hash_init_122_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_121_s0  (
	.D(\top/hash_out [121]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [121])
);
defparam \top/processor/core_hash_init_121_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_120_s0  (
	.D(\top/hash_out [120]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [120])
);
defparam \top/processor/core_hash_init_120_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_119_s0  (
	.D(\top/hash_out [119]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [119])
);
defparam \top/processor/core_hash_init_119_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_118_s0  (
	.D(\top/hash_out [118]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [118])
);
defparam \top/processor/core_hash_init_118_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_117_s0  (
	.D(\top/hash_out [117]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [117])
);
defparam \top/processor/core_hash_init_117_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_116_s0  (
	.D(\top/hash_out [116]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [116])
);
defparam \top/processor/core_hash_init_116_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_115_s0  (
	.D(\top/hash_out [115]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [115])
);
defparam \top/processor/core_hash_init_115_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_114_s0  (
	.D(\top/hash_out [114]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [114])
);
defparam \top/processor/core_hash_init_114_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_113_s0  (
	.D(\top/hash_out [113]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [113])
);
defparam \top/processor/core_hash_init_113_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_112_s0  (
	.D(\top/hash_out [112]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [112])
);
defparam \top/processor/core_hash_init_112_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_111_s0  (
	.D(\top/hash_out [111]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [111])
);
defparam \top/processor/core_hash_init_111_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_110_s0  (
	.D(\top/hash_out [110]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [110])
);
defparam \top/processor/core_hash_init_110_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_109_s0  (
	.D(\top/hash_out [109]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [109])
);
defparam \top/processor/core_hash_init_109_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_108_s0  (
	.D(\top/hash_out [108]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [108])
);
defparam \top/processor/core_hash_init_108_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_107_s0  (
	.D(\top/hash_out [107]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [107])
);
defparam \top/processor/core_hash_init_107_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_106_s0  (
	.D(\top/hash_out [106]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [106])
);
defparam \top/processor/core_hash_init_106_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_105_s0  (
	.D(\top/hash_out [105]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [105])
);
defparam \top/processor/core_hash_init_105_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_104_s0  (
	.D(\top/hash_out [104]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [104])
);
defparam \top/processor/core_hash_init_104_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_103_s0  (
	.D(\top/hash_out [103]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [103])
);
defparam \top/processor/core_hash_init_103_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_102_s0  (
	.D(\top/hash_out [102]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [102])
);
defparam \top/processor/core_hash_init_102_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_101_s0  (
	.D(\top/hash_out [101]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [101])
);
defparam \top/processor/core_hash_init_101_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_100_s0  (
	.D(\top/hash_out [100]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [100])
);
defparam \top/processor/core_hash_init_100_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_99_s0  (
	.D(\top/hash_out [99]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [99])
);
defparam \top/processor/core_hash_init_99_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_98_s0  (
	.D(\top/hash_out [98]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [98])
);
defparam \top/processor/core_hash_init_98_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_97_s0  (
	.D(\top/hash_out [97]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [97])
);
defparam \top/processor/core_hash_init_97_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_96_s0  (
	.D(\top/hash_out [96]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [96])
);
defparam \top/processor/core_hash_init_96_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_95_s0  (
	.D(\top/hash_out [95]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [95])
);
defparam \top/processor/core_hash_init_95_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_94_s0  (
	.D(\top/hash_out [94]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [94])
);
defparam \top/processor/core_hash_init_94_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_93_s0  (
	.D(\top/hash_out [93]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [93])
);
defparam \top/processor/core_hash_init_93_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_92_s0  (
	.D(\top/hash_out [92]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [92])
);
defparam \top/processor/core_hash_init_92_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_91_s0  (
	.D(\top/hash_out [91]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [91])
);
defparam \top/processor/core_hash_init_91_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_90_s0  (
	.D(\top/hash_out [90]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [90])
);
defparam \top/processor/core_hash_init_90_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_89_s0  (
	.D(\top/hash_out [89]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [89])
);
defparam \top/processor/core_hash_init_89_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_88_s0  (
	.D(\top/hash_out [88]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [88])
);
defparam \top/processor/core_hash_init_88_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_87_s0  (
	.D(\top/hash_out [87]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [87])
);
defparam \top/processor/core_hash_init_87_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_86_s0  (
	.D(\top/hash_out [86]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [86])
);
defparam \top/processor/core_hash_init_86_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_85_s0  (
	.D(\top/hash_out [85]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [85])
);
defparam \top/processor/core_hash_init_85_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_84_s0  (
	.D(\top/hash_out [84]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [84])
);
defparam \top/processor/core_hash_init_84_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_83_s0  (
	.D(\top/hash_out [83]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [83])
);
defparam \top/processor/core_hash_init_83_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_82_s0  (
	.D(\top/hash_out [82]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [82])
);
defparam \top/processor/core_hash_init_82_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_81_s0  (
	.D(\top/hash_out [81]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [81])
);
defparam \top/processor/core_hash_init_81_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_80_s0  (
	.D(\top/hash_out [80]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [80])
);
defparam \top/processor/core_hash_init_80_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_79_s0  (
	.D(\top/hash_out [79]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [79])
);
defparam \top/processor/core_hash_init_79_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_78_s0  (
	.D(\top/hash_out [78]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [78])
);
defparam \top/processor/core_hash_init_78_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_77_s0  (
	.D(\top/hash_out [77]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [77])
);
defparam \top/processor/core_hash_init_77_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_76_s0  (
	.D(\top/hash_out [76]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [76])
);
defparam \top/processor/core_hash_init_76_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_75_s0  (
	.D(\top/hash_out [75]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [75])
);
defparam \top/processor/core_hash_init_75_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_74_s0  (
	.D(\top/hash_out [74]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [74])
);
defparam \top/processor/core_hash_init_74_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_73_s0  (
	.D(\top/hash_out [73]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [73])
);
defparam \top/processor/core_hash_init_73_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_72_s0  (
	.D(\top/hash_out [72]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [72])
);
defparam \top/processor/core_hash_init_72_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_71_s0  (
	.D(\top/hash_out [71]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [71])
);
defparam \top/processor/core_hash_init_71_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_70_s0  (
	.D(\top/hash_out [70]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [70])
);
defparam \top/processor/core_hash_init_70_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_69_s0  (
	.D(\top/hash_out [69]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [69])
);
defparam \top/processor/core_hash_init_69_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_68_s0  (
	.D(\top/hash_out [68]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [68])
);
defparam \top/processor/core_hash_init_68_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_67_s0  (
	.D(\top/hash_out [67]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [67])
);
defparam \top/processor/core_hash_init_67_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_66_s0  (
	.D(\top/hash_out [66]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [66])
);
defparam \top/processor/core_hash_init_66_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_65_s0  (
	.D(\top/hash_out [65]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [65])
);
defparam \top/processor/core_hash_init_65_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_64_s0  (
	.D(\top/hash_out [64]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [64])
);
defparam \top/processor/core_hash_init_64_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_63_s0  (
	.D(\top/hash_out [63]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [63])
);
defparam \top/processor/core_hash_init_63_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_62_s0  (
	.D(\top/hash_out [62]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [62])
);
defparam \top/processor/core_hash_init_62_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_61_s0  (
	.D(\top/hash_out [61]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [61])
);
defparam \top/processor/core_hash_init_61_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_60_s0  (
	.D(\top/hash_out [60]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [60])
);
defparam \top/processor/core_hash_init_60_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_59_s0  (
	.D(\top/hash_out [59]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [59])
);
defparam \top/processor/core_hash_init_59_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_58_s0  (
	.D(\top/hash_out [58]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [58])
);
defparam \top/processor/core_hash_init_58_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_57_s0  (
	.D(\top/hash_out [57]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [57])
);
defparam \top/processor/core_hash_init_57_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_56_s0  (
	.D(\top/hash_out [56]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [56])
);
defparam \top/processor/core_hash_init_56_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_55_s0  (
	.D(\top/hash_out [55]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [55])
);
defparam \top/processor/core_hash_init_55_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_54_s0  (
	.D(\top/hash_out [54]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [54])
);
defparam \top/processor/core_hash_init_54_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_53_s0  (
	.D(\top/hash_out [53]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [53])
);
defparam \top/processor/core_hash_init_53_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_52_s0  (
	.D(\top/hash_out [52]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [52])
);
defparam \top/processor/core_hash_init_52_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_51_s0  (
	.D(\top/hash_out [51]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [51])
);
defparam \top/processor/core_hash_init_51_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_50_s0  (
	.D(\top/hash_out [50]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [50])
);
defparam \top/processor/core_hash_init_50_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_49_s0  (
	.D(\top/hash_out [49]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [49])
);
defparam \top/processor/core_hash_init_49_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_48_s0  (
	.D(\top/hash_out [48]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [48])
);
defparam \top/processor/core_hash_init_48_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_47_s0  (
	.D(\top/hash_out [47]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [47])
);
defparam \top/processor/core_hash_init_47_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_46_s0  (
	.D(\top/hash_out [46]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [46])
);
defparam \top/processor/core_hash_init_46_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_45_s0  (
	.D(\top/hash_out [45]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [45])
);
defparam \top/processor/core_hash_init_45_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_44_s0  (
	.D(\top/hash_out [44]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [44])
);
defparam \top/processor/core_hash_init_44_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_43_s0  (
	.D(\top/hash_out [43]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [43])
);
defparam \top/processor/core_hash_init_43_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_42_s0  (
	.D(\top/hash_out [42]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [42])
);
defparam \top/processor/core_hash_init_42_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_41_s0  (
	.D(\top/hash_out [41]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [41])
);
defparam \top/processor/core_hash_init_41_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_40_s0  (
	.D(\top/hash_out [40]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [40])
);
defparam \top/processor/core_hash_init_40_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_39_s0  (
	.D(\top/hash_out [39]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [39])
);
defparam \top/processor/core_hash_init_39_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_38_s0  (
	.D(\top/hash_out [38]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [38])
);
defparam \top/processor/core_hash_init_38_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_37_s0  (
	.D(\top/hash_out [37]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [37])
);
defparam \top/processor/core_hash_init_37_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_36_s0  (
	.D(\top/hash_out [36]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [36])
);
defparam \top/processor/core_hash_init_36_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_35_s0  (
	.D(\top/hash_out [35]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [35])
);
defparam \top/processor/core_hash_init_35_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_34_s0  (
	.D(\top/hash_out [34]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [34])
);
defparam \top/processor/core_hash_init_34_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_33_s0  (
	.D(\top/hash_out [33]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [33])
);
defparam \top/processor/core_hash_init_33_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_32_s0  (
	.D(\top/hash_out [32]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [32])
);
defparam \top/processor/core_hash_init_32_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_31_s0  (
	.D(\top/hash_out [31]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [31])
);
defparam \top/processor/core_hash_init_31_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_30_s0  (
	.D(\top/hash_out [30]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [30])
);
defparam \top/processor/core_hash_init_30_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_29_s0  (
	.D(\top/hash_out [29]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [29])
);
defparam \top/processor/core_hash_init_29_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_28_s0  (
	.D(\top/hash_out [28]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [28])
);
defparam \top/processor/core_hash_init_28_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_27_s0  (
	.D(\top/hash_out [27]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [27])
);
defparam \top/processor/core_hash_init_27_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_26_s0  (
	.D(\top/hash_out [26]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [26])
);
defparam \top/processor/core_hash_init_26_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_25_s0  (
	.D(\top/hash_out [25]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [25])
);
defparam \top/processor/core_hash_init_25_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_24_s0  (
	.D(\top/hash_out [24]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [24])
);
defparam \top/processor/core_hash_init_24_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_23_s0  (
	.D(\top/hash_out [23]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [23])
);
defparam \top/processor/core_hash_init_23_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_22_s0  (
	.D(\top/hash_out [22]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [22])
);
defparam \top/processor/core_hash_init_22_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_21_s0  (
	.D(\top/hash_out [21]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [21])
);
defparam \top/processor/core_hash_init_21_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_20_s0  (
	.D(\top/hash_out [20]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [20])
);
defparam \top/processor/core_hash_init_20_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_19_s0  (
	.D(\top/hash_out [19]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [19])
);
defparam \top/processor/core_hash_init_19_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_18_s0  (
	.D(\top/hash_out [18]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [18])
);
defparam \top/processor/core_hash_init_18_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_17_s0  (
	.D(\top/hash_out [17]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [17])
);
defparam \top/processor/core_hash_init_17_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_16_s0  (
	.D(\top/hash_out [16]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [16])
);
defparam \top/processor/core_hash_init_16_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_15_s0  (
	.D(\top/hash_out [15]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [15])
);
defparam \top/processor/core_hash_init_15_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_14_s0  (
	.D(\top/hash_out [14]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [14])
);
defparam \top/processor/core_hash_init_14_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_13_s0  (
	.D(\top/hash_out [13]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [13])
);
defparam \top/processor/core_hash_init_13_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_12_s0  (
	.D(\top/hash_out [12]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [12])
);
defparam \top/processor/core_hash_init_12_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_11_s0  (
	.D(\top/hash_out [11]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [11])
);
defparam \top/processor/core_hash_init_11_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_10_s0  (
	.D(\top/hash_out [10]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [10])
);
defparam \top/processor/core_hash_init_10_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_9_s0  (
	.D(\top/hash_out [9]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [9])
);
defparam \top/processor/core_hash_init_9_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_8_s0  (
	.D(\top/hash_out [8]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [8])
);
defparam \top/processor/core_hash_init_8_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_7_s0  (
	.D(\top/hash_out [7]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [7])
);
defparam \top/processor/core_hash_init_7_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_6_s0  (
	.D(\top/hash_out [6]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [6])
);
defparam \top/processor/core_hash_init_6_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_5_s0  (
	.D(\top/hash_out [5]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [5])
);
defparam \top/processor/core_hash_init_5_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_4_s0  (
	.D(\top/hash_out [4]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [4])
);
defparam \top/processor/core_hash_init_4_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_3_s0  (
	.D(\top/hash_out [3]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [3])
);
defparam \top/processor/core_hash_init_3_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_2_s0  (
	.D(\top/hash_out [2]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [2])
);
defparam \top/processor/core_hash_init_2_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_1_s0  (
	.D(\top/hash_out [1]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [1])
);
defparam \top/processor/core_hash_init_1_s0 .INIT=1'b0;
DFFCE \top/processor/core_hash_init_0_s0  (
	.D(\top/hash_out [0]),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_init [0])
);
defparam \top/processor/core_hash_init_0_s0 .INIT=1'b0;
DFFCE \top/processor/core_use_init_s0  (
	.D(VCC),
	.CLK(clk),
	.CE(\top/processor/n9790_13 ),
	.CLEAR(rst),
	.Q(\top/processor/core_use_init )
);
defparam \top/processor/core_use_init_s0 .INIT=1'b0;
DFFCE \top/processor/core_busy_s0  (
	.D(\top/processor/n8408_6 ),
	.CLK(clk),
	.CE(\top/processor/core_busy_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_busy )
);
defparam \top/processor/core_busy_s0 .INIT=1'b0;
DFFCE \top/processor/core_ready_prev_s0  (
	.D(\top/processor/core_ready ),
	.CLK(clk),
	.CE(\top/processor/n9790_15 ),
	.CLEAR(rst),
	.Q(\top/processor/core_ready_prev )
);
defparam \top/processor/core_ready_prev_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_255_s0  (
	.D(\top/processor/n10561_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [255])
);
defparam \top/processor/hash_state_255_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_253_s0  (
	.D(\top/processor/n10563_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [253])
);
defparam \top/processor/hash_state_253_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_252_s0  (
	.D(\top/processor/n10564_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [252])
);
defparam \top/processor/hash_state_252_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_251_s0  (
	.D(\top/processor/n10565_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [251])
);
defparam \top/processor/hash_state_251_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_250_s0  (
	.D(\top/processor/n10566_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [250])
);
defparam \top/processor/hash_state_250_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_249_s0  (
	.D(\top/processor/n10567_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [249])
);
defparam \top/processor/hash_state_249_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_248_s0  (
	.D(\top/processor/n10568_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [248])
);
defparam \top/processor/hash_state_248_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_247_s0  (
	.D(\top/processor/n10569_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [247])
);
defparam \top/processor/hash_state_247_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_246_s0  (
	.D(\top/processor/n10570_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [246])
);
defparam \top/processor/hash_state_246_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_245_s0  (
	.D(\top/processor/n10571_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [245])
);
defparam \top/processor/hash_state_245_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_244_s0  (
	.D(\top/processor/n10572_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [244])
);
defparam \top/processor/hash_state_244_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_243_s0  (
	.D(\top/processor/n10573_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [243])
);
defparam \top/processor/hash_state_243_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_242_s0  (
	.D(\top/processor/n10574_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [242])
);
defparam \top/processor/hash_state_242_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_241_s0  (
	.D(\top/processor/n10575_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [241])
);
defparam \top/processor/hash_state_241_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_240_s0  (
	.D(\top/processor/n10576_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [240])
);
defparam \top/processor/hash_state_240_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_239_s0  (
	.D(\top/processor/n10577_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [239])
);
defparam \top/processor/hash_state_239_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_238_s0  (
	.D(\top/processor/n10578_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [238])
);
defparam \top/processor/hash_state_238_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_237_s0  (
	.D(\top/processor/n10579_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [237])
);
defparam \top/processor/hash_state_237_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_236_s0  (
	.D(\top/processor/n10580_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [236])
);
defparam \top/processor/hash_state_236_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_235_s0  (
	.D(\top/processor/n10581_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [235])
);
defparam \top/processor/hash_state_235_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_234_s0  (
	.D(\top/processor/n10582_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [234])
);
defparam \top/processor/hash_state_234_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_233_s0  (
	.D(\top/processor/n10583_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [233])
);
defparam \top/processor/hash_state_233_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_232_s0  (
	.D(\top/processor/n10584_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [232])
);
defparam \top/processor/hash_state_232_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_231_s0  (
	.D(\top/processor/n10585_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [231])
);
defparam \top/processor/hash_state_231_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_230_s0  (
	.D(\top/processor/n10586_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [230])
);
defparam \top/processor/hash_state_230_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_229_s0  (
	.D(\top/processor/n10587_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [229])
);
defparam \top/processor/hash_state_229_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_228_s0  (
	.D(\top/processor/n10588_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [228])
);
defparam \top/processor/hash_state_228_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_227_s0  (
	.D(\top/processor/n10589_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [227])
);
defparam \top/processor/hash_state_227_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_226_s0  (
	.D(\top/processor/n10590_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [226])
);
defparam \top/processor/hash_state_226_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_225_s0  (
	.D(\top/processor/n10591_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [225])
);
defparam \top/processor/hash_state_225_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_224_s0  (
	.D(\top/processor/n10592_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [224])
);
defparam \top/processor/hash_state_224_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_223_s0  (
	.D(\top/processor/n10593_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [223])
);
defparam \top/processor/hash_state_223_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_222_s0  (
	.D(\top/processor/n10594_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [222])
);
defparam \top/processor/hash_state_222_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_221_s0  (
	.D(\top/processor/n10595_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [221])
);
defparam \top/processor/hash_state_221_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_220_s0  (
	.D(\top/processor/n10596_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [220])
);
defparam \top/processor/hash_state_220_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_219_s0  (
	.D(\top/processor/n10597_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [219])
);
defparam \top/processor/hash_state_219_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_218_s0  (
	.D(\top/processor/n10598_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [218])
);
defparam \top/processor/hash_state_218_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_217_s0  (
	.D(\top/processor/n10599_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [217])
);
defparam \top/processor/hash_state_217_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_216_s0  (
	.D(\top/processor/n10600_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [216])
);
defparam \top/processor/hash_state_216_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_215_s0  (
	.D(\top/processor/n10601_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [215])
);
defparam \top/processor/hash_state_215_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_214_s0  (
	.D(\top/processor/n10602_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [214])
);
defparam \top/processor/hash_state_214_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_213_s0  (
	.D(\top/processor/n10603_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [213])
);
defparam \top/processor/hash_state_213_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_212_s0  (
	.D(\top/processor/n10604_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [212])
);
defparam \top/processor/hash_state_212_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_211_s0  (
	.D(\top/processor/n10605_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [211])
);
defparam \top/processor/hash_state_211_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_210_s0  (
	.D(\top/processor/n10606_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [210])
);
defparam \top/processor/hash_state_210_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_209_s0  (
	.D(\top/processor/n10607_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [209])
);
defparam \top/processor/hash_state_209_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_208_s0  (
	.D(\top/processor/n10608_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [208])
);
defparam \top/processor/hash_state_208_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_207_s0  (
	.D(\top/processor/n10609_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [207])
);
defparam \top/processor/hash_state_207_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_206_s0  (
	.D(\top/processor/n10610_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [206])
);
defparam \top/processor/hash_state_206_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_205_s0  (
	.D(\top/processor/n10611_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [205])
);
defparam \top/processor/hash_state_205_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_204_s0  (
	.D(\top/processor/n10612_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [204])
);
defparam \top/processor/hash_state_204_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_203_s0  (
	.D(\top/processor/n10613_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [203])
);
defparam \top/processor/hash_state_203_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_202_s0  (
	.D(\top/processor/n10614_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [202])
);
defparam \top/processor/hash_state_202_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_201_s0  (
	.D(\top/processor/n10615_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [201])
);
defparam \top/processor/hash_state_201_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_200_s0  (
	.D(\top/processor/n10616_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [200])
);
defparam \top/processor/hash_state_200_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_199_s0  (
	.D(\top/processor/n10617_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [199])
);
defparam \top/processor/hash_state_199_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_198_s0  (
	.D(\top/processor/n10618_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [198])
);
defparam \top/processor/hash_state_198_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_197_s0  (
	.D(\top/processor/n10619_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [197])
);
defparam \top/processor/hash_state_197_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_196_s0  (
	.D(\top/processor/n10620_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [196])
);
defparam \top/processor/hash_state_196_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_195_s0  (
	.D(\top/processor/n10621_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [195])
);
defparam \top/processor/hash_state_195_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_194_s0  (
	.D(\top/processor/n10622_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [194])
);
defparam \top/processor/hash_state_194_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_193_s0  (
	.D(\top/processor/n10623_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [193])
);
defparam \top/processor/hash_state_193_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_192_s0  (
	.D(\top/processor/n10624_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [192])
);
defparam \top/processor/hash_state_192_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_191_s0  (
	.D(\top/processor/n10625_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [191])
);
defparam \top/processor/hash_state_191_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_190_s0  (
	.D(\top/processor/n10626_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [190])
);
defparam \top/processor/hash_state_190_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_189_s0  (
	.D(\top/processor/n10627_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [189])
);
defparam \top/processor/hash_state_189_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_188_s0  (
	.D(\top/processor/n10628_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [188])
);
defparam \top/processor/hash_state_188_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_187_s0  (
	.D(\top/processor/n10629_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [187])
);
defparam \top/processor/hash_state_187_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_186_s0  (
	.D(\top/processor/n10630_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [186])
);
defparam \top/processor/hash_state_186_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_185_s0  (
	.D(\top/processor/n10631_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [185])
);
defparam \top/processor/hash_state_185_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_184_s0  (
	.D(\top/processor/n10632_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [184])
);
defparam \top/processor/hash_state_184_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_183_s0  (
	.D(\top/processor/n10633_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [183])
);
defparam \top/processor/hash_state_183_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_182_s0  (
	.D(\top/processor/n10634_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [182])
);
defparam \top/processor/hash_state_182_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_181_s0  (
	.D(\top/processor/n10635_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [181])
);
defparam \top/processor/hash_state_181_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_180_s0  (
	.D(\top/processor/n10636_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [180])
);
defparam \top/processor/hash_state_180_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_179_s0  (
	.D(\top/processor/n10637_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [179])
);
defparam \top/processor/hash_state_179_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_178_s0  (
	.D(\top/processor/n10638_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [178])
);
defparam \top/processor/hash_state_178_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_177_s0  (
	.D(\top/processor/n10639_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [177])
);
defparam \top/processor/hash_state_177_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_176_s0  (
	.D(\top/processor/n10640_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [176])
);
defparam \top/processor/hash_state_176_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_175_s0  (
	.D(\top/processor/n10641_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [175])
);
defparam \top/processor/hash_state_175_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_174_s0  (
	.D(\top/processor/n10642_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [174])
);
defparam \top/processor/hash_state_174_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_173_s0  (
	.D(\top/processor/n10643_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [173])
);
defparam \top/processor/hash_state_173_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_172_s0  (
	.D(\top/processor/n10644_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [172])
);
defparam \top/processor/hash_state_172_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_171_s0  (
	.D(\top/processor/n10645_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [171])
);
defparam \top/processor/hash_state_171_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_170_s0  (
	.D(\top/processor/n10646_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [170])
);
defparam \top/processor/hash_state_170_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_169_s0  (
	.D(\top/processor/n10647_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [169])
);
defparam \top/processor/hash_state_169_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_168_s0  (
	.D(\top/processor/n10648_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [168])
);
defparam \top/processor/hash_state_168_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_167_s0  (
	.D(\top/processor/n10649_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [167])
);
defparam \top/processor/hash_state_167_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_166_s0  (
	.D(\top/processor/n10650_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [166])
);
defparam \top/processor/hash_state_166_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_165_s0  (
	.D(\top/processor/n10651_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [165])
);
defparam \top/processor/hash_state_165_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_164_s0  (
	.D(\top/processor/n10652_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [164])
);
defparam \top/processor/hash_state_164_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_163_s0  (
	.D(\top/processor/n10653_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [163])
);
defparam \top/processor/hash_state_163_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_162_s0  (
	.D(\top/processor/n10654_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [162])
);
defparam \top/processor/hash_state_162_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_161_s0  (
	.D(\top/processor/n10655_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [161])
);
defparam \top/processor/hash_state_161_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_160_s0  (
	.D(\top/processor/n10656_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [160])
);
defparam \top/processor/hash_state_160_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_159_s0  (
	.D(\top/processor/n10657_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [159])
);
defparam \top/processor/hash_state_159_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_158_s0  (
	.D(\top/processor/n10658_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [158])
);
defparam \top/processor/hash_state_158_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_157_s0  (
	.D(\top/processor/n10659_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [157])
);
defparam \top/processor/hash_state_157_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_156_s0  (
	.D(\top/processor/n10660_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [156])
);
defparam \top/processor/hash_state_156_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_155_s0  (
	.D(\top/processor/n10661_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [155])
);
defparam \top/processor/hash_state_155_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_154_s0  (
	.D(\top/processor/n10662_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [154])
);
defparam \top/processor/hash_state_154_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_153_s0  (
	.D(\top/processor/n10663_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [153])
);
defparam \top/processor/hash_state_153_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_152_s0  (
	.D(\top/processor/n10664_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [152])
);
defparam \top/processor/hash_state_152_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_151_s0  (
	.D(\top/processor/n10665_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [151])
);
defparam \top/processor/hash_state_151_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_150_s0  (
	.D(\top/processor/n10666_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [150])
);
defparam \top/processor/hash_state_150_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_149_s0  (
	.D(\top/processor/n10667_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [149])
);
defparam \top/processor/hash_state_149_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_148_s0  (
	.D(\top/processor/n10668_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [148])
);
defparam \top/processor/hash_state_148_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_147_s0  (
	.D(\top/processor/n10669_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [147])
);
defparam \top/processor/hash_state_147_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_146_s0  (
	.D(\top/processor/n10670_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [146])
);
defparam \top/processor/hash_state_146_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_145_s0  (
	.D(\top/processor/n10671_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [145])
);
defparam \top/processor/hash_state_145_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_144_s0  (
	.D(\top/processor/n10672_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [144])
);
defparam \top/processor/hash_state_144_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_143_s0  (
	.D(\top/processor/n10673_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [143])
);
defparam \top/processor/hash_state_143_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_142_s0  (
	.D(\top/processor/n10674_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [142])
);
defparam \top/processor/hash_state_142_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_141_s0  (
	.D(\top/processor/n10675_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [141])
);
defparam \top/processor/hash_state_141_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_140_s0  (
	.D(\top/processor/n10676_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [140])
);
defparam \top/processor/hash_state_140_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_139_s0  (
	.D(\top/processor/n10677_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [139])
);
defparam \top/processor/hash_state_139_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_138_s0  (
	.D(\top/processor/n10678_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [138])
);
defparam \top/processor/hash_state_138_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_137_s0  (
	.D(\top/processor/n10679_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [137])
);
defparam \top/processor/hash_state_137_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_136_s0  (
	.D(\top/processor/n10680_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [136])
);
defparam \top/processor/hash_state_136_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_135_s0  (
	.D(\top/processor/n10681_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [135])
);
defparam \top/processor/hash_state_135_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_134_s0  (
	.D(\top/processor/n10682_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [134])
);
defparam \top/processor/hash_state_134_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_133_s0  (
	.D(\top/processor/n10683_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [133])
);
defparam \top/processor/hash_state_133_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_132_s0  (
	.D(\top/processor/n10684_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [132])
);
defparam \top/processor/hash_state_132_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_131_s0  (
	.D(\top/processor/n10685_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [131])
);
defparam \top/processor/hash_state_131_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_130_s0  (
	.D(\top/processor/n10686_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [130])
);
defparam \top/processor/hash_state_130_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_129_s0  (
	.D(\top/processor/n10687_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [129])
);
defparam \top/processor/hash_state_129_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_128_s0  (
	.D(\top/processor/n10688_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [128])
);
defparam \top/processor/hash_state_128_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_127_s0  (
	.D(\top/processor/n10689_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [127])
);
defparam \top/processor/hash_state_127_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_126_s0  (
	.D(\top/processor/n10690_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [126])
);
defparam \top/processor/hash_state_126_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_125_s0  (
	.D(\top/processor/n10691_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [125])
);
defparam \top/processor/hash_state_125_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_124_s0  (
	.D(\top/processor/n10692_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [124])
);
defparam \top/processor/hash_state_124_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_123_s0  (
	.D(\top/processor/n10693_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [123])
);
defparam \top/processor/hash_state_123_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_122_s0  (
	.D(\top/processor/n10694_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [122])
);
defparam \top/processor/hash_state_122_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_121_s0  (
	.D(\top/processor/n10695_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [121])
);
defparam \top/processor/hash_state_121_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_120_s0  (
	.D(\top/processor/n10696_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [120])
);
defparam \top/processor/hash_state_120_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_119_s0  (
	.D(\top/processor/n10697_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [119])
);
defparam \top/processor/hash_state_119_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_118_s0  (
	.D(\top/processor/n10698_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [118])
);
defparam \top/processor/hash_state_118_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_117_s0  (
	.D(\top/processor/n10699_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [117])
);
defparam \top/processor/hash_state_117_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_116_s0  (
	.D(\top/processor/n10700_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [116])
);
defparam \top/processor/hash_state_116_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_115_s0  (
	.D(\top/processor/n10701_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [115])
);
defparam \top/processor/hash_state_115_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_114_s0  (
	.D(\top/processor/n10702_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [114])
);
defparam \top/processor/hash_state_114_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_113_s0  (
	.D(\top/processor/n10703_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [113])
);
defparam \top/processor/hash_state_113_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_112_s0  (
	.D(\top/processor/n10704_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [112])
);
defparam \top/processor/hash_state_112_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_111_s0  (
	.D(\top/processor/n10705_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [111])
);
defparam \top/processor/hash_state_111_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_110_s0  (
	.D(\top/processor/n10706_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [110])
);
defparam \top/processor/hash_state_110_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_109_s0  (
	.D(\top/processor/n10707_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [109])
);
defparam \top/processor/hash_state_109_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_108_s0  (
	.D(\top/processor/n10708_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [108])
);
defparam \top/processor/hash_state_108_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_107_s0  (
	.D(\top/processor/n10709_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [107])
);
defparam \top/processor/hash_state_107_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_106_s0  (
	.D(\top/processor/n10710_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [106])
);
defparam \top/processor/hash_state_106_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_105_s0  (
	.D(\top/processor/n10711_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [105])
);
defparam \top/processor/hash_state_105_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_104_s0  (
	.D(\top/processor/n10712_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [104])
);
defparam \top/processor/hash_state_104_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_103_s0  (
	.D(\top/processor/n10713_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [103])
);
defparam \top/processor/hash_state_103_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_102_s0  (
	.D(\top/processor/n10714_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [102])
);
defparam \top/processor/hash_state_102_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_101_s0  (
	.D(\top/processor/n10715_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [101])
);
defparam \top/processor/hash_state_101_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_100_s0  (
	.D(\top/processor/n10716_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [100])
);
defparam \top/processor/hash_state_100_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_99_s0  (
	.D(\top/processor/n10717_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [99])
);
defparam \top/processor/hash_state_99_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_98_s0  (
	.D(\top/processor/n10718_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [98])
);
defparam \top/processor/hash_state_98_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_97_s0  (
	.D(\top/processor/n10719_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [97])
);
defparam \top/processor/hash_state_97_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_96_s0  (
	.D(\top/processor/n10720_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [96])
);
defparam \top/processor/hash_state_96_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_95_s0  (
	.D(\top/processor/n10721_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [95])
);
defparam \top/processor/hash_state_95_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_94_s0  (
	.D(\top/processor/n10722_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [94])
);
defparam \top/processor/hash_state_94_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_93_s0  (
	.D(\top/processor/n10723_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [93])
);
defparam \top/processor/hash_state_93_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_92_s0  (
	.D(\top/processor/n10724_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [92])
);
defparam \top/processor/hash_state_92_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_91_s0  (
	.D(\top/processor/n10725_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [91])
);
defparam \top/processor/hash_state_91_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_90_s0  (
	.D(\top/processor/n10726_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [90])
);
defparam \top/processor/hash_state_90_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_89_s0  (
	.D(\top/processor/n10727_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [89])
);
defparam \top/processor/hash_state_89_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_88_s0  (
	.D(\top/processor/n10728_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [88])
);
defparam \top/processor/hash_state_88_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_87_s0  (
	.D(\top/processor/n10729_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [87])
);
defparam \top/processor/hash_state_87_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_86_s0  (
	.D(\top/processor/n10730_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [86])
);
defparam \top/processor/hash_state_86_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_85_s0  (
	.D(\top/processor/n10731_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [85])
);
defparam \top/processor/hash_state_85_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_84_s0  (
	.D(\top/processor/n10732_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [84])
);
defparam \top/processor/hash_state_84_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_83_s0  (
	.D(\top/processor/n10733_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [83])
);
defparam \top/processor/hash_state_83_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_82_s0  (
	.D(\top/processor/n10734_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [82])
);
defparam \top/processor/hash_state_82_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_81_s0  (
	.D(\top/processor/n10735_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [81])
);
defparam \top/processor/hash_state_81_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_80_s0  (
	.D(\top/processor/n10736_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [80])
);
defparam \top/processor/hash_state_80_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_79_s0  (
	.D(\top/processor/n10737_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [79])
);
defparam \top/processor/hash_state_79_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_78_s0  (
	.D(\top/processor/n10738_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [78])
);
defparam \top/processor/hash_state_78_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_77_s0  (
	.D(\top/processor/n10739_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [77])
);
defparam \top/processor/hash_state_77_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_76_s0  (
	.D(\top/processor/n10740_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [76])
);
defparam \top/processor/hash_state_76_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_75_s0  (
	.D(\top/processor/n10741_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [75])
);
defparam \top/processor/hash_state_75_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_74_s0  (
	.D(\top/processor/n10742_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [74])
);
defparam \top/processor/hash_state_74_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_73_s0  (
	.D(\top/processor/n10743_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [73])
);
defparam \top/processor/hash_state_73_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_72_s0  (
	.D(\top/processor/n10744_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [72])
);
defparam \top/processor/hash_state_72_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_71_s0  (
	.D(\top/processor/n10745_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [71])
);
defparam \top/processor/hash_state_71_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_70_s0  (
	.D(\top/processor/n10746_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [70])
);
defparam \top/processor/hash_state_70_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_69_s0  (
	.D(\top/processor/n10747_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [69])
);
defparam \top/processor/hash_state_69_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_68_s0  (
	.D(\top/processor/n10748_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [68])
);
defparam \top/processor/hash_state_68_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_67_s0  (
	.D(\top/processor/n10749_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [67])
);
defparam \top/processor/hash_state_67_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_66_s0  (
	.D(\top/processor/n10750_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [66])
);
defparam \top/processor/hash_state_66_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_65_s0  (
	.D(\top/processor/n10751_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [65])
);
defparam \top/processor/hash_state_65_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_64_s0  (
	.D(\top/processor/n10752_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [64])
);
defparam \top/processor/hash_state_64_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_63_s0  (
	.D(\top/processor/n10753_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [63])
);
defparam \top/processor/hash_state_63_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_62_s0  (
	.D(\top/processor/n10754_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [62])
);
defparam \top/processor/hash_state_62_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_61_s0  (
	.D(\top/processor/n10755_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [61])
);
defparam \top/processor/hash_state_61_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_60_s0  (
	.D(\top/processor/n10756_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [60])
);
defparam \top/processor/hash_state_60_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_59_s0  (
	.D(\top/processor/n10757_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [59])
);
defparam \top/processor/hash_state_59_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_58_s0  (
	.D(\top/processor/n10758_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [58])
);
defparam \top/processor/hash_state_58_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_57_s0  (
	.D(\top/processor/n10759_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [57])
);
defparam \top/processor/hash_state_57_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_56_s0  (
	.D(\top/processor/n10760_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [56])
);
defparam \top/processor/hash_state_56_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_55_s0  (
	.D(\top/processor/n10761_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [55])
);
defparam \top/processor/hash_state_55_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_54_s0  (
	.D(\top/processor/n10762_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [54])
);
defparam \top/processor/hash_state_54_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_53_s0  (
	.D(\top/processor/n10763_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [53])
);
defparam \top/processor/hash_state_53_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_52_s0  (
	.D(\top/processor/n10764_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [52])
);
defparam \top/processor/hash_state_52_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_51_s0  (
	.D(\top/processor/n10765_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [51])
);
defparam \top/processor/hash_state_51_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_50_s0  (
	.D(\top/processor/n10766_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [50])
);
defparam \top/processor/hash_state_50_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_49_s0  (
	.D(\top/processor/n10767_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [49])
);
defparam \top/processor/hash_state_49_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_48_s0  (
	.D(\top/processor/n10768_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [48])
);
defparam \top/processor/hash_state_48_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_47_s0  (
	.D(\top/processor/n10769_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [47])
);
defparam \top/processor/hash_state_47_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_46_s0  (
	.D(\top/processor/n10770_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [46])
);
defparam \top/processor/hash_state_46_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_45_s0  (
	.D(\top/processor/n10771_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [45])
);
defparam \top/processor/hash_state_45_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_44_s0  (
	.D(\top/processor/n10772_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [44])
);
defparam \top/processor/hash_state_44_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_43_s0  (
	.D(\top/processor/n10773_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [43])
);
defparam \top/processor/hash_state_43_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_42_s0  (
	.D(\top/processor/n10774_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [42])
);
defparam \top/processor/hash_state_42_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_41_s0  (
	.D(\top/processor/n10775_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [41])
);
defparam \top/processor/hash_state_41_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_40_s0  (
	.D(\top/processor/n10776_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [40])
);
defparam \top/processor/hash_state_40_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_39_s0  (
	.D(\top/processor/n10777_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [39])
);
defparam \top/processor/hash_state_39_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_38_s0  (
	.D(\top/processor/n10778_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [38])
);
defparam \top/processor/hash_state_38_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_37_s0  (
	.D(\top/processor/n10779_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [37])
);
defparam \top/processor/hash_state_37_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_36_s0  (
	.D(\top/processor/n10780_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [36])
);
defparam \top/processor/hash_state_36_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_35_s0  (
	.D(\top/processor/n10781_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [35])
);
defparam \top/processor/hash_state_35_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_34_s0  (
	.D(\top/processor/n10782_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [34])
);
defparam \top/processor/hash_state_34_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_33_s0  (
	.D(\top/processor/n10783_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [33])
);
defparam \top/processor/hash_state_33_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_32_s0  (
	.D(\top/processor/n10784_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [32])
);
defparam \top/processor/hash_state_32_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_31_s0  (
	.D(\top/processor/n10785_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [31])
);
defparam \top/processor/hash_state_31_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_30_s0  (
	.D(\top/processor/n10786_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [30])
);
defparam \top/processor/hash_state_30_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_29_s0  (
	.D(\top/processor/n10787_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [29])
);
defparam \top/processor/hash_state_29_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_28_s0  (
	.D(\top/processor/n10788_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [28])
);
defparam \top/processor/hash_state_28_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_27_s0  (
	.D(\top/processor/n10789_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [27])
);
defparam \top/processor/hash_state_27_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_26_s0  (
	.D(\top/processor/n10790_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [26])
);
defparam \top/processor/hash_state_26_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_25_s0  (
	.D(\top/processor/n10791_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [25])
);
defparam \top/processor/hash_state_25_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_24_s0  (
	.D(\top/processor/n10792_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [24])
);
defparam \top/processor/hash_state_24_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_23_s0  (
	.D(\top/processor/n10793_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [23])
);
defparam \top/processor/hash_state_23_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_22_s0  (
	.D(\top/processor/n10794_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [22])
);
defparam \top/processor/hash_state_22_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_21_s0  (
	.D(\top/processor/n10795_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [21])
);
defparam \top/processor/hash_state_21_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_20_s0  (
	.D(\top/processor/n10796_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [20])
);
defparam \top/processor/hash_state_20_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_19_s0  (
	.D(\top/processor/n10797_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [19])
);
defparam \top/processor/hash_state_19_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_18_s0  (
	.D(\top/processor/n10798_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [18])
);
defparam \top/processor/hash_state_18_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_17_s0  (
	.D(\top/processor/n10799_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [17])
);
defparam \top/processor/hash_state_17_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_16_s0  (
	.D(\top/processor/n10800_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [16])
);
defparam \top/processor/hash_state_16_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_15_s0  (
	.D(\top/processor/n10801_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [15])
);
defparam \top/processor/hash_state_15_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_14_s0  (
	.D(\top/processor/n10802_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [14])
);
defparam \top/processor/hash_state_14_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_13_s0  (
	.D(\top/processor/n10803_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [13])
);
defparam \top/processor/hash_state_13_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_12_s0  (
	.D(\top/processor/n10804_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [12])
);
defparam \top/processor/hash_state_12_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_11_s0  (
	.D(\top/processor/n10805_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [11])
);
defparam \top/processor/hash_state_11_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_10_s0  (
	.D(\top/processor/n10806_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [10])
);
defparam \top/processor/hash_state_10_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_9_s0  (
	.D(\top/processor/n10807_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [9])
);
defparam \top/processor/hash_state_9_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_8_s0  (
	.D(\top/processor/n10808_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [8])
);
defparam \top/processor/hash_state_8_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_7_s0  (
	.D(\top/processor/n10809_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [7])
);
defparam \top/processor/hash_state_7_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_6_s0  (
	.D(\top/processor/n10810_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [6])
);
defparam \top/processor/hash_state_6_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_5_s0  (
	.D(\top/processor/n10811_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [5])
);
defparam \top/processor/hash_state_5_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_4_s0  (
	.D(\top/processor/n10812_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [4])
);
defparam \top/processor/hash_state_4_s0 .INIT=1'b1;
DFFPE \top/processor/hash_state_3_s0  (
	.D(\top/processor/n10813_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [3])
);
defparam \top/processor/hash_state_3_s0 .INIT=1'b1;
DFFCE \top/processor/hash_state_2_s0  (
	.D(\top/processor/n10814_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [2])
);
defparam \top/processor/hash_state_2_s0 .INIT=1'b0;
DFFCE \top/processor/hash_state_1_s0  (
	.D(\top/processor/n10815_15 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.CLEAR(rst),
	.Q(\top/hash_out [1])
);
defparam \top/processor/hash_state_1_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_0_s0  (
	.D(\top/processor/n10816_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [0])
);
defparam \top/processor/hash_state_0_s0 .INIT=1'b1;
DFFCE \top/processor/total_bits_63_s0  (
	.D(\top/processor/n11378_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [63])
);
defparam \top/processor/total_bits_63_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_62_s0  (
	.D(\top/processor/n11379_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [62])
);
defparam \top/processor/total_bits_62_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_61_s0  (
	.D(\top/processor/n11380_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [61])
);
defparam \top/processor/total_bits_61_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_60_s0  (
	.D(\top/processor/n11381_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [60])
);
defparam \top/processor/total_bits_60_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_59_s0  (
	.D(\top/processor/n11382_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [59])
);
defparam \top/processor/total_bits_59_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_58_s0  (
	.D(\top/processor/n11383_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [58])
);
defparam \top/processor/total_bits_58_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_57_s0  (
	.D(\top/processor/n11384_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [57])
);
defparam \top/processor/total_bits_57_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_56_s0  (
	.D(\top/processor/n11385_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [56])
);
defparam \top/processor/total_bits_56_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_55_s0  (
	.D(\top/processor/n11386_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [55])
);
defparam \top/processor/total_bits_55_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_54_s0  (
	.D(\top/processor/n11387_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [54])
);
defparam \top/processor/total_bits_54_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_53_s0  (
	.D(\top/processor/n11388_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [53])
);
defparam \top/processor/total_bits_53_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_52_s0  (
	.D(\top/processor/n11389_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [52])
);
defparam \top/processor/total_bits_52_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_51_s0  (
	.D(\top/processor/n11390_18 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [51])
);
defparam \top/processor/total_bits_51_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_50_s0  (
	.D(\top/processor/n11391_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [50])
);
defparam \top/processor/total_bits_50_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_49_s0  (
	.D(\top/processor/n11392_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [49])
);
defparam \top/processor/total_bits_49_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_48_s0  (
	.D(\top/processor/n11393_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [48])
);
defparam \top/processor/total_bits_48_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_47_s0  (
	.D(\top/processor/n11394_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [47])
);
defparam \top/processor/total_bits_47_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_46_s0  (
	.D(\top/processor/n11395_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [46])
);
defparam \top/processor/total_bits_46_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_45_s0  (
	.D(\top/processor/n11396_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [45])
);
defparam \top/processor/total_bits_45_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_44_s0  (
	.D(\top/processor/n11397_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [44])
);
defparam \top/processor/total_bits_44_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_43_s0  (
	.D(\top/processor/n11398_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [43])
);
defparam \top/processor/total_bits_43_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_42_s0  (
	.D(\top/processor/n11399_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [42])
);
defparam \top/processor/total_bits_42_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_41_s0  (
	.D(\top/processor/n11400_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [41])
);
defparam \top/processor/total_bits_41_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_40_s0  (
	.D(\top/processor/n11401_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [40])
);
defparam \top/processor/total_bits_40_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_39_s0  (
	.D(\top/processor/n11402_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [39])
);
defparam \top/processor/total_bits_39_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_38_s0  (
	.D(\top/processor/n11403_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [38])
);
defparam \top/processor/total_bits_38_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_37_s0  (
	.D(\top/processor/n11404_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [37])
);
defparam \top/processor/total_bits_37_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_36_s0  (
	.D(\top/processor/n11405_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [36])
);
defparam \top/processor/total_bits_36_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_35_s0  (
	.D(\top/processor/n11406_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [35])
);
defparam \top/processor/total_bits_35_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_34_s0  (
	.D(\top/processor/n11407_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [34])
);
defparam \top/processor/total_bits_34_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_33_s0  (
	.D(\top/processor/n11408_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [33])
);
defparam \top/processor/total_bits_33_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_32_s0  (
	.D(\top/processor/n11409_17 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [32])
);
defparam \top/processor/total_bits_32_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_31_s0  (
	.D(\top/processor/n11410_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [31])
);
defparam \top/processor/total_bits_31_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_30_s0  (
	.D(\top/processor/n11411_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [30])
);
defparam \top/processor/total_bits_30_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_29_s0  (
	.D(\top/processor/n11412_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [29])
);
defparam \top/processor/total_bits_29_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_28_s0  (
	.D(\top/processor/n11413_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [28])
);
defparam \top/processor/total_bits_28_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_27_s0  (
	.D(\top/processor/n11414_17 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [27])
);
defparam \top/processor/total_bits_27_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_26_s0  (
	.D(\top/processor/n11415_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [26])
);
defparam \top/processor/total_bits_26_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_25_s0  (
	.D(\top/processor/n11416_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [25])
);
defparam \top/processor/total_bits_25_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_24_s0  (
	.D(\top/processor/n11417_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [24])
);
defparam \top/processor/total_bits_24_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_23_s0  (
	.D(\top/processor/n11418_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [23])
);
defparam \top/processor/total_bits_23_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_22_s0  (
	.D(\top/processor/n11419_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [22])
);
defparam \top/processor/total_bits_22_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_21_s0  (
	.D(\top/processor/n11420_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [21])
);
defparam \top/processor/total_bits_21_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_20_s0  (
	.D(\top/processor/n11421_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [20])
);
defparam \top/processor/total_bits_20_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_19_s0  (
	.D(\top/processor/n11422_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [19])
);
defparam \top/processor/total_bits_19_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_18_s0  (
	.D(\top/processor/n11423_17 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [18])
);
defparam \top/processor/total_bits_18_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_17_s0  (
	.D(\top/processor/n11424_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [17])
);
defparam \top/processor/total_bits_17_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_16_s0  (
	.D(\top/processor/n11425_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [16])
);
defparam \top/processor/total_bits_16_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_15_s0  (
	.D(\top/processor/n11426_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [15])
);
defparam \top/processor/total_bits_15_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_14_s0  (
	.D(\top/processor/n11427_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [14])
);
defparam \top/processor/total_bits_14_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_13_s0  (
	.D(\top/processor/n11428_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [13])
);
defparam \top/processor/total_bits_13_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_12_s0  (
	.D(\top/processor/n11429_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [12])
);
defparam \top/processor/total_bits_12_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_11_s0  (
	.D(\top/processor/n11430_17 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [11])
);
defparam \top/processor/total_bits_11_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_10_s0  (
	.D(\top/processor/n11431_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [10])
);
defparam \top/processor/total_bits_10_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_9_s0  (
	.D(\top/processor/n11432_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [9])
);
defparam \top/processor/total_bits_9_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_8_s0  (
	.D(\top/processor/n11433_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [8])
);
defparam \top/processor/total_bits_8_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_7_s0  (
	.D(\top/processor/n11434_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [7])
);
defparam \top/processor/total_bits_7_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_6_s0  (
	.D(\top/processor/n11435_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [6])
);
defparam \top/processor/total_bits_6_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_5_s0  (
	.D(\top/processor/n11436_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [5])
);
defparam \top/processor/total_bits_5_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_4_s0  (
	.D(\top/processor/n11437_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [4])
);
defparam \top/processor/total_bits_4_s0 .INIT=1'b0;
DFFCE \top/processor/total_bits_3_s0  (
	.D(\top/processor/n11438_14 ),
	.CLK(clk),
	.CE(\top/processor/total_bits_63_8 ),
	.CLEAR(rst),
	.Q(\top/processor/total_bits [3])
);
defparam \top/processor/total_bits_3_s0 .INIT=1'b0;
DFFCE \top/processor/seen_last_s0  (
	.D(\top/state_0 [0]),
	.CLK(clk),
	.CE(\top/processor/seen_last_8 ),
	.CLEAR(rst),
	.Q(\top/processor/seen_last )
);
defparam \top/processor/seen_last_s0 .INIT=1'b0;
DFFCE \top/processor/need_length_block_s0  (
	.D(\top/processor/n11361_16 ),
	.CLK(clk),
	.CE(\top/processor/need_length_block_8 ),
	.CLEAR(rst),
	.Q(\top/processor/need_length_block )
);
defparam \top/processor/need_length_block_s0 .INIT=1'b0;
DFFCE \top/processor/pad_index_5_s0  (
	.D(\top/processor/n11372_14 ),
	.CLK(clk),
	.CE(\top/processor/pad_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/pad_index [5])
);
defparam \top/processor/pad_index_5_s0 .INIT=1'b0;
DFFCE \top/processor/pad_index_4_s0  (
	.D(\top/processor/n11373_14 ),
	.CLK(clk),
	.CE(\top/processor/pad_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/pad_index [4])
);
defparam \top/processor/pad_index_4_s0 .INIT=1'b0;
DFFCE \top/processor/pad_index_3_s0  (
	.D(\top/processor/n11374_14 ),
	.CLK(clk),
	.CE(\top/processor/pad_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/pad_index [3])
);
defparam \top/processor/pad_index_3_s0 .INIT=1'b0;
DFFCE \top/processor/pad_index_2_s0  (
	.D(\top/processor/n11375_14 ),
	.CLK(clk),
	.CE(\top/processor/pad_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/pad_index [2])
);
defparam \top/processor/pad_index_2_s0 .INIT=1'b0;
DFFCE \top/processor/pad_index_1_s0  (
	.D(\top/processor/n11376_14 ),
	.CLK(clk),
	.CE(\top/processor/pad_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/pad_index [1])
);
defparam \top/processor/pad_index_1_s0 .INIT=1'b0;
DFFCE \top/processor/pad_index_0_s0  (
	.D(\top/processor/n11377_14 ),
	.CLK(clk),
	.CE(\top/processor/pad_index_5_8 ),
	.CLEAR(rst),
	.Q(\top/processor/pad_index [0])
);
defparam \top/processor/pad_index_0_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_511_s0  (
	.D(\top/processor/n10817_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [511])
);
defparam \top/processor/block_buffer_511_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_510_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [510])
);
defparam \top/processor/block_buffer_510_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_509_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [509])
);
defparam \top/processor/block_buffer_509_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_508_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [508])
);
defparam \top/processor/block_buffer_508_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_507_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [507])
);
defparam \top/processor/block_buffer_507_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_506_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [506])
);
defparam \top/processor/block_buffer_506_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_505_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [505])
);
defparam \top/processor/block_buffer_505_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_504_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_511_15 ),
	.Q(\top/processor/block_buffer [504])
);
defparam \top/processor/block_buffer_504_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_503_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [503])
);
defparam \top/processor/block_buffer_503_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_502_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [502])
);
defparam \top/processor/block_buffer_502_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_501_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [501])
);
defparam \top/processor/block_buffer_501_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_500_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [500])
);
defparam \top/processor/block_buffer_500_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_499_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [499])
);
defparam \top/processor/block_buffer_499_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_498_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [498])
);
defparam \top/processor/block_buffer_498_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_497_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [497])
);
defparam \top/processor/block_buffer_497_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_496_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_503_8 ),
	.Q(\top/processor/block_buffer [496])
);
defparam \top/processor/block_buffer_496_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_495_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [495])
);
defparam \top/processor/block_buffer_495_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_494_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [494])
);
defparam \top/processor/block_buffer_494_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_493_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [493])
);
defparam \top/processor/block_buffer_493_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_492_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [492])
);
defparam \top/processor/block_buffer_492_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_491_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [491])
);
defparam \top/processor/block_buffer_491_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_490_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [490])
);
defparam \top/processor/block_buffer_490_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_489_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [489])
);
defparam \top/processor/block_buffer_489_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_488_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_495_8 ),
	.Q(\top/processor/block_buffer [488])
);
defparam \top/processor/block_buffer_488_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_487_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [487])
);
defparam \top/processor/block_buffer_487_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_486_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [486])
);
defparam \top/processor/block_buffer_486_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_485_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [485])
);
defparam \top/processor/block_buffer_485_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_484_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [484])
);
defparam \top/processor/block_buffer_484_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_483_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [483])
);
defparam \top/processor/block_buffer_483_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_482_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [482])
);
defparam \top/processor/block_buffer_482_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_481_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [481])
);
defparam \top/processor/block_buffer_481_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_480_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_487_8 ),
	.Q(\top/processor/block_buffer [480])
);
defparam \top/processor/block_buffer_480_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_479_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [479])
);
defparam \top/processor/block_buffer_479_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_478_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [478])
);
defparam \top/processor/block_buffer_478_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_477_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [477])
);
defparam \top/processor/block_buffer_477_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_476_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [476])
);
defparam \top/processor/block_buffer_476_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_475_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [475])
);
defparam \top/processor/block_buffer_475_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_474_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [474])
);
defparam \top/processor/block_buffer_474_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_473_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [473])
);
defparam \top/processor/block_buffer_473_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_472_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_479_8 ),
	.Q(\top/processor/block_buffer [472])
);
defparam \top/processor/block_buffer_472_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_471_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [471])
);
defparam \top/processor/block_buffer_471_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_470_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [470])
);
defparam \top/processor/block_buffer_470_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_469_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [469])
);
defparam \top/processor/block_buffer_469_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_468_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [468])
);
defparam \top/processor/block_buffer_468_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_467_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [467])
);
defparam \top/processor/block_buffer_467_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_466_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [466])
);
defparam \top/processor/block_buffer_466_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_465_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [465])
);
defparam \top/processor/block_buffer_465_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_464_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_471_8 ),
	.Q(\top/processor/block_buffer [464])
);
defparam \top/processor/block_buffer_464_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_463_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [463])
);
defparam \top/processor/block_buffer_463_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_462_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [462])
);
defparam \top/processor/block_buffer_462_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_461_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [461])
);
defparam \top/processor/block_buffer_461_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_460_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [460])
);
defparam \top/processor/block_buffer_460_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_459_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [459])
);
defparam \top/processor/block_buffer_459_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_458_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [458])
);
defparam \top/processor/block_buffer_458_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_457_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [457])
);
defparam \top/processor/block_buffer_457_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_456_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_463_8 ),
	.Q(\top/processor/block_buffer [456])
);
defparam \top/processor/block_buffer_456_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_455_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [455])
);
defparam \top/processor/block_buffer_455_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_454_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [454])
);
defparam \top/processor/block_buffer_454_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_453_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [453])
);
defparam \top/processor/block_buffer_453_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_452_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [452])
);
defparam \top/processor/block_buffer_452_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_451_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [451])
);
defparam \top/processor/block_buffer_451_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_450_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [450])
);
defparam \top/processor/block_buffer_450_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_449_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [449])
);
defparam \top/processor/block_buffer_449_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_448_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_455_8 ),
	.Q(\top/processor/block_buffer [448])
);
defparam \top/processor/block_buffer_448_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_447_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [447])
);
defparam \top/processor/block_buffer_447_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_446_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [446])
);
defparam \top/processor/block_buffer_446_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_445_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [445])
);
defparam \top/processor/block_buffer_445_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_444_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [444])
);
defparam \top/processor/block_buffer_444_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_443_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [443])
);
defparam \top/processor/block_buffer_443_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_442_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [442])
);
defparam \top/processor/block_buffer_442_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_441_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [441])
);
defparam \top/processor/block_buffer_441_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_440_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_447_14 ),
	.Q(\top/processor/block_buffer [440])
);
defparam \top/processor/block_buffer_440_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_439_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [439])
);
defparam \top/processor/block_buffer_439_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_438_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [438])
);
defparam \top/processor/block_buffer_438_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_437_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [437])
);
defparam \top/processor/block_buffer_437_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_436_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [436])
);
defparam \top/processor/block_buffer_436_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_435_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [435])
);
defparam \top/processor/block_buffer_435_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_434_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [434])
);
defparam \top/processor/block_buffer_434_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_433_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [433])
);
defparam \top/processor/block_buffer_433_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_432_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_439_8 ),
	.Q(\top/processor/block_buffer [432])
);
defparam \top/processor/block_buffer_432_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_431_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [431])
);
defparam \top/processor/block_buffer_431_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_430_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [430])
);
defparam \top/processor/block_buffer_430_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_429_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [429])
);
defparam \top/processor/block_buffer_429_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_428_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [428])
);
defparam \top/processor/block_buffer_428_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_427_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [427])
);
defparam \top/processor/block_buffer_427_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_426_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [426])
);
defparam \top/processor/block_buffer_426_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_425_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [425])
);
defparam \top/processor/block_buffer_425_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_424_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_431_8 ),
	.Q(\top/processor/block_buffer [424])
);
defparam \top/processor/block_buffer_424_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_423_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [423])
);
defparam \top/processor/block_buffer_423_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_422_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [422])
);
defparam \top/processor/block_buffer_422_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_421_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [421])
);
defparam \top/processor/block_buffer_421_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_420_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [420])
);
defparam \top/processor/block_buffer_420_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_419_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [419])
);
defparam \top/processor/block_buffer_419_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_418_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [418])
);
defparam \top/processor/block_buffer_418_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_417_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [417])
);
defparam \top/processor/block_buffer_417_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_416_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_423_8 ),
	.Q(\top/processor/block_buffer [416])
);
defparam \top/processor/block_buffer_416_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_415_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [415])
);
defparam \top/processor/block_buffer_415_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_414_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [414])
);
defparam \top/processor/block_buffer_414_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_413_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [413])
);
defparam \top/processor/block_buffer_413_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_412_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [412])
);
defparam \top/processor/block_buffer_412_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_411_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [411])
);
defparam \top/processor/block_buffer_411_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_410_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [410])
);
defparam \top/processor/block_buffer_410_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_409_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [409])
);
defparam \top/processor/block_buffer_409_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_408_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_415_8 ),
	.Q(\top/processor/block_buffer [408])
);
defparam \top/processor/block_buffer_408_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_407_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [407])
);
defparam \top/processor/block_buffer_407_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_406_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [406])
);
defparam \top/processor/block_buffer_406_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_405_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [405])
);
defparam \top/processor/block_buffer_405_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_404_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [404])
);
defparam \top/processor/block_buffer_404_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_403_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [403])
);
defparam \top/processor/block_buffer_403_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_402_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [402])
);
defparam \top/processor/block_buffer_402_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_401_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [401])
);
defparam \top/processor/block_buffer_401_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_400_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_407_8 ),
	.Q(\top/processor/block_buffer [400])
);
defparam \top/processor/block_buffer_400_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_399_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [399])
);
defparam \top/processor/block_buffer_399_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_398_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [398])
);
defparam \top/processor/block_buffer_398_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_397_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [397])
);
defparam \top/processor/block_buffer_397_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_396_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [396])
);
defparam \top/processor/block_buffer_396_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_395_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [395])
);
defparam \top/processor/block_buffer_395_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_394_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [394])
);
defparam \top/processor/block_buffer_394_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_393_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [393])
);
defparam \top/processor/block_buffer_393_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_392_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_399_8 ),
	.Q(\top/processor/block_buffer [392])
);
defparam \top/processor/block_buffer_392_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_391_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [391])
);
defparam \top/processor/block_buffer_391_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_390_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [390])
);
defparam \top/processor/block_buffer_390_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_389_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [389])
);
defparam \top/processor/block_buffer_389_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_388_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [388])
);
defparam \top/processor/block_buffer_388_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_387_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [387])
);
defparam \top/processor/block_buffer_387_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_386_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [386])
);
defparam \top/processor/block_buffer_386_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_385_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [385])
);
defparam \top/processor/block_buffer_385_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_384_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_391_8 ),
	.Q(\top/processor/block_buffer [384])
);
defparam \top/processor/block_buffer_384_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_383_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [383])
);
defparam \top/processor/block_buffer_383_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_382_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [382])
);
defparam \top/processor/block_buffer_382_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_381_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [381])
);
defparam \top/processor/block_buffer_381_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_380_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [380])
);
defparam \top/processor/block_buffer_380_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_379_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [379])
);
defparam \top/processor/block_buffer_379_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_378_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [378])
);
defparam \top/processor/block_buffer_378_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_377_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [377])
);
defparam \top/processor/block_buffer_377_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_376_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_383_13 ),
	.Q(\top/processor/block_buffer [376])
);
defparam \top/processor/block_buffer_376_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_375_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [375])
);
defparam \top/processor/block_buffer_375_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_374_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [374])
);
defparam \top/processor/block_buffer_374_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_373_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [373])
);
defparam \top/processor/block_buffer_373_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_372_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [372])
);
defparam \top/processor/block_buffer_372_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_371_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [371])
);
defparam \top/processor/block_buffer_371_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_370_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [370])
);
defparam \top/processor/block_buffer_370_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_369_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [369])
);
defparam \top/processor/block_buffer_369_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_368_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_375_8 ),
	.Q(\top/processor/block_buffer [368])
);
defparam \top/processor/block_buffer_368_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_367_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [367])
);
defparam \top/processor/block_buffer_367_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_366_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [366])
);
defparam \top/processor/block_buffer_366_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_365_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [365])
);
defparam \top/processor/block_buffer_365_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_364_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [364])
);
defparam \top/processor/block_buffer_364_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_363_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [363])
);
defparam \top/processor/block_buffer_363_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_362_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [362])
);
defparam \top/processor/block_buffer_362_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_361_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [361])
);
defparam \top/processor/block_buffer_361_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_360_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_367_8 ),
	.Q(\top/processor/block_buffer [360])
);
defparam \top/processor/block_buffer_360_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_359_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [359])
);
defparam \top/processor/block_buffer_359_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_358_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [358])
);
defparam \top/processor/block_buffer_358_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_357_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [357])
);
defparam \top/processor/block_buffer_357_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_356_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [356])
);
defparam \top/processor/block_buffer_356_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_355_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [355])
);
defparam \top/processor/block_buffer_355_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_354_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [354])
);
defparam \top/processor/block_buffer_354_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_353_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [353])
);
defparam \top/processor/block_buffer_353_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_352_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_359_8 ),
	.Q(\top/processor/block_buffer [352])
);
defparam \top/processor/block_buffer_352_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_351_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [351])
);
defparam \top/processor/block_buffer_351_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_350_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [350])
);
defparam \top/processor/block_buffer_350_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_349_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [349])
);
defparam \top/processor/block_buffer_349_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_348_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [348])
);
defparam \top/processor/block_buffer_348_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_347_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [347])
);
defparam \top/processor/block_buffer_347_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_346_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [346])
);
defparam \top/processor/block_buffer_346_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_345_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [345])
);
defparam \top/processor/block_buffer_345_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_344_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_351_8 ),
	.Q(\top/processor/block_buffer [344])
);
defparam \top/processor/block_buffer_344_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_343_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [343])
);
defparam \top/processor/block_buffer_343_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_342_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [342])
);
defparam \top/processor/block_buffer_342_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_341_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [341])
);
defparam \top/processor/block_buffer_341_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_340_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [340])
);
defparam \top/processor/block_buffer_340_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_339_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [339])
);
defparam \top/processor/block_buffer_339_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_338_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [338])
);
defparam \top/processor/block_buffer_338_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_337_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [337])
);
defparam \top/processor/block_buffer_337_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_336_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_343_8 ),
	.Q(\top/processor/block_buffer [336])
);
defparam \top/processor/block_buffer_336_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_335_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [335])
);
defparam \top/processor/block_buffer_335_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_334_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [334])
);
defparam \top/processor/block_buffer_334_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_333_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [333])
);
defparam \top/processor/block_buffer_333_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_332_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [332])
);
defparam \top/processor/block_buffer_332_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_331_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [331])
);
defparam \top/processor/block_buffer_331_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_330_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [330])
);
defparam \top/processor/block_buffer_330_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_329_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [329])
);
defparam \top/processor/block_buffer_329_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_328_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_335_8 ),
	.Q(\top/processor/block_buffer [328])
);
defparam \top/processor/block_buffer_328_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_327_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [327])
);
defparam \top/processor/block_buffer_327_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_326_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [326])
);
defparam \top/processor/block_buffer_326_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_325_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [325])
);
defparam \top/processor/block_buffer_325_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_324_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [324])
);
defparam \top/processor/block_buffer_324_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_323_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [323])
);
defparam \top/processor/block_buffer_323_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_322_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [322])
);
defparam \top/processor/block_buffer_322_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_321_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [321])
);
defparam \top/processor/block_buffer_321_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_320_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_327_8 ),
	.Q(\top/processor/block_buffer [320])
);
defparam \top/processor/block_buffer_320_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_319_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [319])
);
defparam \top/processor/block_buffer_319_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_318_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [318])
);
defparam \top/processor/block_buffer_318_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_317_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [317])
);
defparam \top/processor/block_buffer_317_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_316_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [316])
);
defparam \top/processor/block_buffer_316_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_315_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [315])
);
defparam \top/processor/block_buffer_315_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_314_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [314])
);
defparam \top/processor/block_buffer_314_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_313_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [313])
);
defparam \top/processor/block_buffer_313_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_312_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_319_8 ),
	.Q(\top/processor/block_buffer [312])
);
defparam \top/processor/block_buffer_312_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_311_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [311])
);
defparam \top/processor/block_buffer_311_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_310_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [310])
);
defparam \top/processor/block_buffer_310_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_309_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [309])
);
defparam \top/processor/block_buffer_309_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_308_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [308])
);
defparam \top/processor/block_buffer_308_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_307_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [307])
);
defparam \top/processor/block_buffer_307_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_306_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [306])
);
defparam \top/processor/block_buffer_306_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_305_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [305])
);
defparam \top/processor/block_buffer_305_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_304_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_311_8 ),
	.Q(\top/processor/block_buffer [304])
);
defparam \top/processor/block_buffer_304_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_303_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [303])
);
defparam \top/processor/block_buffer_303_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_302_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [302])
);
defparam \top/processor/block_buffer_302_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_301_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [301])
);
defparam \top/processor/block_buffer_301_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_300_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [300])
);
defparam \top/processor/block_buffer_300_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_299_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [299])
);
defparam \top/processor/block_buffer_299_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_298_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [298])
);
defparam \top/processor/block_buffer_298_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_297_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [297])
);
defparam \top/processor/block_buffer_297_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_296_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_303_8 ),
	.Q(\top/processor/block_buffer [296])
);
defparam \top/processor/block_buffer_296_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_295_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [295])
);
defparam \top/processor/block_buffer_295_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_294_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [294])
);
defparam \top/processor/block_buffer_294_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_293_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [293])
);
defparam \top/processor/block_buffer_293_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_292_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [292])
);
defparam \top/processor/block_buffer_292_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_291_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [291])
);
defparam \top/processor/block_buffer_291_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_290_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [290])
);
defparam \top/processor/block_buffer_290_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_289_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [289])
);
defparam \top/processor/block_buffer_289_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_288_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_295_8 ),
	.Q(\top/processor/block_buffer [288])
);
defparam \top/processor/block_buffer_288_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_287_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [287])
);
defparam \top/processor/block_buffer_287_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_286_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [286])
);
defparam \top/processor/block_buffer_286_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_285_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [285])
);
defparam \top/processor/block_buffer_285_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_284_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [284])
);
defparam \top/processor/block_buffer_284_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_283_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [283])
);
defparam \top/processor/block_buffer_283_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_282_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [282])
);
defparam \top/processor/block_buffer_282_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_281_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [281])
);
defparam \top/processor/block_buffer_281_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_280_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_287_8 ),
	.Q(\top/processor/block_buffer [280])
);
defparam \top/processor/block_buffer_280_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_279_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [279])
);
defparam \top/processor/block_buffer_279_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_278_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [278])
);
defparam \top/processor/block_buffer_278_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_277_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [277])
);
defparam \top/processor/block_buffer_277_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_276_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [276])
);
defparam \top/processor/block_buffer_276_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_275_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [275])
);
defparam \top/processor/block_buffer_275_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_274_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [274])
);
defparam \top/processor/block_buffer_274_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_273_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [273])
);
defparam \top/processor/block_buffer_273_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_272_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_279_8 ),
	.Q(\top/processor/block_buffer [272])
);
defparam \top/processor/block_buffer_272_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_271_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [271])
);
defparam \top/processor/block_buffer_271_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_270_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [270])
);
defparam \top/processor/block_buffer_270_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_269_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [269])
);
defparam \top/processor/block_buffer_269_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_268_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [268])
);
defparam \top/processor/block_buffer_268_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_267_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [267])
);
defparam \top/processor/block_buffer_267_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_266_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [266])
);
defparam \top/processor/block_buffer_266_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_265_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [265])
);
defparam \top/processor/block_buffer_265_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_264_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_271_8 ),
	.Q(\top/processor/block_buffer [264])
);
defparam \top/processor/block_buffer_264_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_263_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [263])
);
defparam \top/processor/block_buffer_263_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_262_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [262])
);
defparam \top/processor/block_buffer_262_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_261_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [261])
);
defparam \top/processor/block_buffer_261_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_260_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [260])
);
defparam \top/processor/block_buffer_260_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_259_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [259])
);
defparam \top/processor/block_buffer_259_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_258_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [258])
);
defparam \top/processor/block_buffer_258_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_257_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [257])
);
defparam \top/processor/block_buffer_257_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_256_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_263_8 ),
	.Q(\top/processor/block_buffer [256])
);
defparam \top/processor/block_buffer_256_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_255_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [255])
);
defparam \top/processor/block_buffer_255_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_254_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [254])
);
defparam \top/processor/block_buffer_254_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_253_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [253])
);
defparam \top/processor/block_buffer_253_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_252_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [252])
);
defparam \top/processor/block_buffer_252_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_251_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [251])
);
defparam \top/processor/block_buffer_251_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_250_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [250])
);
defparam \top/processor/block_buffer_250_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_249_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [249])
);
defparam \top/processor/block_buffer_249_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_248_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_255_13 ),
	.Q(\top/processor/block_buffer [248])
);
defparam \top/processor/block_buffer_248_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_247_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [247])
);
defparam \top/processor/block_buffer_247_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_246_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [246])
);
defparam \top/processor/block_buffer_246_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_245_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [245])
);
defparam \top/processor/block_buffer_245_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_244_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [244])
);
defparam \top/processor/block_buffer_244_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_243_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [243])
);
defparam \top/processor/block_buffer_243_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_242_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [242])
);
defparam \top/processor/block_buffer_242_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_241_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [241])
);
defparam \top/processor/block_buffer_241_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_240_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_247_8 ),
	.Q(\top/processor/block_buffer [240])
);
defparam \top/processor/block_buffer_240_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_239_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [239])
);
defparam \top/processor/block_buffer_239_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_238_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [238])
);
defparam \top/processor/block_buffer_238_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_237_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [237])
);
defparam \top/processor/block_buffer_237_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_236_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [236])
);
defparam \top/processor/block_buffer_236_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_235_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [235])
);
defparam \top/processor/block_buffer_235_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_234_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [234])
);
defparam \top/processor/block_buffer_234_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_233_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [233])
);
defparam \top/processor/block_buffer_233_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_232_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_239_8 ),
	.Q(\top/processor/block_buffer [232])
);
defparam \top/processor/block_buffer_232_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_231_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [231])
);
defparam \top/processor/block_buffer_231_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_230_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [230])
);
defparam \top/processor/block_buffer_230_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_229_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [229])
);
defparam \top/processor/block_buffer_229_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_228_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [228])
);
defparam \top/processor/block_buffer_228_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_227_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [227])
);
defparam \top/processor/block_buffer_227_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_226_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [226])
);
defparam \top/processor/block_buffer_226_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_225_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [225])
);
defparam \top/processor/block_buffer_225_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_224_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_231_8 ),
	.Q(\top/processor/block_buffer [224])
);
defparam \top/processor/block_buffer_224_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_223_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [223])
);
defparam \top/processor/block_buffer_223_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_222_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [222])
);
defparam \top/processor/block_buffer_222_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_221_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [221])
);
defparam \top/processor/block_buffer_221_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_220_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [220])
);
defparam \top/processor/block_buffer_220_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_219_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [219])
);
defparam \top/processor/block_buffer_219_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_218_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [218])
);
defparam \top/processor/block_buffer_218_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_217_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [217])
);
defparam \top/processor/block_buffer_217_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_216_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_223_8 ),
	.Q(\top/processor/block_buffer [216])
);
defparam \top/processor/block_buffer_216_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_215_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [215])
);
defparam \top/processor/block_buffer_215_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_214_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [214])
);
defparam \top/processor/block_buffer_214_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_213_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [213])
);
defparam \top/processor/block_buffer_213_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_212_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [212])
);
defparam \top/processor/block_buffer_212_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_211_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [211])
);
defparam \top/processor/block_buffer_211_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_210_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [210])
);
defparam \top/processor/block_buffer_210_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_209_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [209])
);
defparam \top/processor/block_buffer_209_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_208_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_215_8 ),
	.Q(\top/processor/block_buffer [208])
);
defparam \top/processor/block_buffer_208_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_207_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [207])
);
defparam \top/processor/block_buffer_207_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_206_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [206])
);
defparam \top/processor/block_buffer_206_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_205_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [205])
);
defparam \top/processor/block_buffer_205_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_204_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [204])
);
defparam \top/processor/block_buffer_204_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_203_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [203])
);
defparam \top/processor/block_buffer_203_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_202_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [202])
);
defparam \top/processor/block_buffer_202_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_201_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [201])
);
defparam \top/processor/block_buffer_201_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_200_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_207_8 ),
	.Q(\top/processor/block_buffer [200])
);
defparam \top/processor/block_buffer_200_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_199_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [199])
);
defparam \top/processor/block_buffer_199_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_198_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [198])
);
defparam \top/processor/block_buffer_198_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_197_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [197])
);
defparam \top/processor/block_buffer_197_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_196_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [196])
);
defparam \top/processor/block_buffer_196_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_195_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [195])
);
defparam \top/processor/block_buffer_195_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_194_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [194])
);
defparam \top/processor/block_buffer_194_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_193_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [193])
);
defparam \top/processor/block_buffer_193_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_192_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_199_8 ),
	.Q(\top/processor/block_buffer [192])
);
defparam \top/processor/block_buffer_192_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_191_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [191])
);
defparam \top/processor/block_buffer_191_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_190_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [190])
);
defparam \top/processor/block_buffer_190_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_189_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [189])
);
defparam \top/processor/block_buffer_189_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_188_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [188])
);
defparam \top/processor/block_buffer_188_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_187_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [187])
);
defparam \top/processor/block_buffer_187_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_186_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [186])
);
defparam \top/processor/block_buffer_186_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_185_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [185])
);
defparam \top/processor/block_buffer_185_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_184_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_191_8 ),
	.Q(\top/processor/block_buffer [184])
);
defparam \top/processor/block_buffer_184_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_183_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [183])
);
defparam \top/processor/block_buffer_183_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_182_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [182])
);
defparam \top/processor/block_buffer_182_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_181_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [181])
);
defparam \top/processor/block_buffer_181_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_180_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [180])
);
defparam \top/processor/block_buffer_180_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_179_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [179])
);
defparam \top/processor/block_buffer_179_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_178_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [178])
);
defparam \top/processor/block_buffer_178_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_177_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [177])
);
defparam \top/processor/block_buffer_177_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_176_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_183_8 ),
	.Q(\top/processor/block_buffer [176])
);
defparam \top/processor/block_buffer_176_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_175_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [175])
);
defparam \top/processor/block_buffer_175_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_174_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [174])
);
defparam \top/processor/block_buffer_174_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_173_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [173])
);
defparam \top/processor/block_buffer_173_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_172_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [172])
);
defparam \top/processor/block_buffer_172_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_171_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [171])
);
defparam \top/processor/block_buffer_171_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_170_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [170])
);
defparam \top/processor/block_buffer_170_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_169_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [169])
);
defparam \top/processor/block_buffer_169_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_168_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_175_8 ),
	.Q(\top/processor/block_buffer [168])
);
defparam \top/processor/block_buffer_168_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_167_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [167])
);
defparam \top/processor/block_buffer_167_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_166_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [166])
);
defparam \top/processor/block_buffer_166_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_165_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [165])
);
defparam \top/processor/block_buffer_165_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_164_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [164])
);
defparam \top/processor/block_buffer_164_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_163_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [163])
);
defparam \top/processor/block_buffer_163_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_162_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [162])
);
defparam \top/processor/block_buffer_162_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_161_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [161])
);
defparam \top/processor/block_buffer_161_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_160_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_167_8 ),
	.Q(\top/processor/block_buffer [160])
);
defparam \top/processor/block_buffer_160_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_159_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [159])
);
defparam \top/processor/block_buffer_159_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_158_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [158])
);
defparam \top/processor/block_buffer_158_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_157_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [157])
);
defparam \top/processor/block_buffer_157_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_156_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [156])
);
defparam \top/processor/block_buffer_156_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_155_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [155])
);
defparam \top/processor/block_buffer_155_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_154_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [154])
);
defparam \top/processor/block_buffer_154_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_153_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [153])
);
defparam \top/processor/block_buffer_153_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_152_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_159_8 ),
	.Q(\top/processor/block_buffer [152])
);
defparam \top/processor/block_buffer_152_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_151_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [151])
);
defparam \top/processor/block_buffer_151_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_150_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [150])
);
defparam \top/processor/block_buffer_150_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_149_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [149])
);
defparam \top/processor/block_buffer_149_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_148_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [148])
);
defparam \top/processor/block_buffer_148_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_147_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [147])
);
defparam \top/processor/block_buffer_147_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_146_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [146])
);
defparam \top/processor/block_buffer_146_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_145_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [145])
);
defparam \top/processor/block_buffer_145_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_144_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_151_8 ),
	.Q(\top/processor/block_buffer [144])
);
defparam \top/processor/block_buffer_144_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_143_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [143])
);
defparam \top/processor/block_buffer_143_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_142_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [142])
);
defparam \top/processor/block_buffer_142_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_141_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [141])
);
defparam \top/processor/block_buffer_141_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_140_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [140])
);
defparam \top/processor/block_buffer_140_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_139_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [139])
);
defparam \top/processor/block_buffer_139_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_138_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [138])
);
defparam \top/processor/block_buffer_138_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_137_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [137])
);
defparam \top/processor/block_buffer_137_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_136_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_143_8 ),
	.Q(\top/processor/block_buffer [136])
);
defparam \top/processor/block_buffer_136_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_135_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [135])
);
defparam \top/processor/block_buffer_135_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_134_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [134])
);
defparam \top/processor/block_buffer_134_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_133_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [133])
);
defparam \top/processor/block_buffer_133_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_132_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [132])
);
defparam \top/processor/block_buffer_132_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_131_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [131])
);
defparam \top/processor/block_buffer_131_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_130_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [130])
);
defparam \top/processor/block_buffer_130_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_129_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [129])
);
defparam \top/processor/block_buffer_129_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_128_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_135_8 ),
	.Q(\top/processor/block_buffer [128])
);
defparam \top/processor/block_buffer_128_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_127_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [127])
);
defparam \top/processor/block_buffer_127_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_126_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [126])
);
defparam \top/processor/block_buffer_126_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_125_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [125])
);
defparam \top/processor/block_buffer_125_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_124_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [124])
);
defparam \top/processor/block_buffer_124_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_123_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [123])
);
defparam \top/processor/block_buffer_123_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_122_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [122])
);
defparam \top/processor/block_buffer_122_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_121_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [121])
);
defparam \top/processor/block_buffer_121_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_120_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_127_8 ),
	.Q(\top/processor/block_buffer [120])
);
defparam \top/processor/block_buffer_120_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_119_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [119])
);
defparam \top/processor/block_buffer_119_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_118_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [118])
);
defparam \top/processor/block_buffer_118_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_117_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [117])
);
defparam \top/processor/block_buffer_117_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_116_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [116])
);
defparam \top/processor/block_buffer_116_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_115_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [115])
);
defparam \top/processor/block_buffer_115_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_114_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [114])
);
defparam \top/processor/block_buffer_114_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_113_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [113])
);
defparam \top/processor/block_buffer_113_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_112_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_119_8 ),
	.Q(\top/processor/block_buffer [112])
);
defparam \top/processor/block_buffer_112_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_111_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [111])
);
defparam \top/processor/block_buffer_111_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_110_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [110])
);
defparam \top/processor/block_buffer_110_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_109_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [109])
);
defparam \top/processor/block_buffer_109_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_108_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [108])
);
defparam \top/processor/block_buffer_108_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_107_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [107])
);
defparam \top/processor/block_buffer_107_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_106_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [106])
);
defparam \top/processor/block_buffer_106_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_105_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [105])
);
defparam \top/processor/block_buffer_105_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_104_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_111_8 ),
	.Q(\top/processor/block_buffer [104])
);
defparam \top/processor/block_buffer_104_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_103_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [103])
);
defparam \top/processor/block_buffer_103_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_102_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [102])
);
defparam \top/processor/block_buffer_102_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_101_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [101])
);
defparam \top/processor/block_buffer_101_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_100_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [100])
);
defparam \top/processor/block_buffer_100_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_99_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [99])
);
defparam \top/processor/block_buffer_99_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_98_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [98])
);
defparam \top/processor/block_buffer_98_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_97_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [97])
);
defparam \top/processor/block_buffer_97_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_96_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_103_8 ),
	.Q(\top/processor/block_buffer [96])
);
defparam \top/processor/block_buffer_96_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_95_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [95])
);
defparam \top/processor/block_buffer_95_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_94_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [94])
);
defparam \top/processor/block_buffer_94_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_93_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [93])
);
defparam \top/processor/block_buffer_93_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_92_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [92])
);
defparam \top/processor/block_buffer_92_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_91_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [91])
);
defparam \top/processor/block_buffer_91_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_90_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [90])
);
defparam \top/processor/block_buffer_90_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_89_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [89])
);
defparam \top/processor/block_buffer_89_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_88_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_95_8 ),
	.Q(\top/processor/block_buffer [88])
);
defparam \top/processor/block_buffer_88_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_87_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [87])
);
defparam \top/processor/block_buffer_87_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_86_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [86])
);
defparam \top/processor/block_buffer_86_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_85_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [85])
);
defparam \top/processor/block_buffer_85_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_84_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [84])
);
defparam \top/processor/block_buffer_84_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_83_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [83])
);
defparam \top/processor/block_buffer_83_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_82_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [82])
);
defparam \top/processor/block_buffer_82_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_81_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [81])
);
defparam \top/processor/block_buffer_81_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_80_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_87_8 ),
	.Q(\top/processor/block_buffer [80])
);
defparam \top/processor/block_buffer_80_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_79_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [79])
);
defparam \top/processor/block_buffer_79_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_78_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [78])
);
defparam \top/processor/block_buffer_78_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_77_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [77])
);
defparam \top/processor/block_buffer_77_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_76_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [76])
);
defparam \top/processor/block_buffer_76_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_75_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [75])
);
defparam \top/processor/block_buffer_75_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_74_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [74])
);
defparam \top/processor/block_buffer_74_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_73_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [73])
);
defparam \top/processor/block_buffer_73_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_72_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_79_8 ),
	.Q(\top/processor/block_buffer [72])
);
defparam \top/processor/block_buffer_72_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_71_s0  (
	.D(\top/processor/n10825_14 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [71])
);
defparam \top/processor/block_buffer_71_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_70_s0  (
	.D(\top/processor/n10818_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [70])
);
defparam \top/processor/block_buffer_70_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_69_s0  (
	.D(\top/processor/n10819_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [69])
);
defparam \top/processor/block_buffer_69_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_68_s0  (
	.D(\top/processor/n10820_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [68])
);
defparam \top/processor/block_buffer_68_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_67_s0  (
	.D(\top/processor/n10821_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [67])
);
defparam \top/processor/block_buffer_67_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_66_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [66])
);
defparam \top/processor/block_buffer_66_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_65_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [65])
);
defparam \top/processor/block_buffer_65_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_64_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_71_8 ),
	.Q(\top/processor/block_buffer [64])
);
defparam \top/processor/block_buffer_64_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_63_s0  (
	.D(\top/processor/n11265_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [63])
);
defparam \top/processor/block_buffer_63_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_62_s0  (
	.D(\top/processor/n11266_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [62])
);
defparam \top/processor/block_buffer_62_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_61_s0  (
	.D(\top/processor/n11267_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [61])
);
defparam \top/processor/block_buffer_61_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_60_s0  (
	.D(\top/processor/n11268_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [60])
);
defparam \top/processor/block_buffer_60_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_59_s0  (
	.D(\top/processor/n11269_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [59])
);
defparam \top/processor/block_buffer_59_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_58_s0  (
	.D(\top/processor/n11270_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [58])
);
defparam \top/processor/block_buffer_58_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_57_s0  (
	.D(\top/processor/n11271_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [57])
);
defparam \top/processor/block_buffer_57_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_56_s0  (
	.D(\top/processor/n11272_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_63_8 ),
	.Q(\top/processor/block_buffer [56])
);
defparam \top/processor/block_buffer_56_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_55_s0  (
	.D(\top/processor/n11273_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [55])
);
defparam \top/processor/block_buffer_55_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_54_s0  (
	.D(\top/processor/n11274_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [54])
);
defparam \top/processor/block_buffer_54_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_53_s0  (
	.D(\top/processor/n11275_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [53])
);
defparam \top/processor/block_buffer_53_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_52_s0  (
	.D(\top/processor/n11276_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [52])
);
defparam \top/processor/block_buffer_52_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_51_s0  (
	.D(\top/processor/n11277_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [51])
);
defparam \top/processor/block_buffer_51_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_50_s0  (
	.D(\top/processor/n11278_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [50])
);
defparam \top/processor/block_buffer_50_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_49_s0  (
	.D(\top/processor/n11279_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [49])
);
defparam \top/processor/block_buffer_49_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_48_s0  (
	.D(\top/processor/n11280_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_55_8 ),
	.Q(\top/processor/block_buffer [48])
);
defparam \top/processor/block_buffer_48_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_47_s0  (
	.D(\top/processor/n11281_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [47])
);
defparam \top/processor/block_buffer_47_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_46_s0  (
	.D(\top/processor/n11282_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [46])
);
defparam \top/processor/block_buffer_46_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_45_s0  (
	.D(\top/processor/n11283_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [45])
);
defparam \top/processor/block_buffer_45_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_44_s0  (
	.D(\top/processor/n11284_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [44])
);
defparam \top/processor/block_buffer_44_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_43_s0  (
	.D(\top/processor/n11285_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [43])
);
defparam \top/processor/block_buffer_43_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_42_s0  (
	.D(\top/processor/n11286_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [42])
);
defparam \top/processor/block_buffer_42_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_41_s0  (
	.D(\top/processor/n11287_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [41])
);
defparam \top/processor/block_buffer_41_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_40_s0  (
	.D(\top/processor/n11288_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_47_8 ),
	.Q(\top/processor/block_buffer [40])
);
defparam \top/processor/block_buffer_40_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_39_s0  (
	.D(\top/processor/n11289_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [39])
);
defparam \top/processor/block_buffer_39_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_38_s0  (
	.D(\top/processor/n11290_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [38])
);
defparam \top/processor/block_buffer_38_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_37_s0  (
	.D(\top/processor/n11291_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [37])
);
defparam \top/processor/block_buffer_37_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_36_s0  (
	.D(\top/processor/n11292_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [36])
);
defparam \top/processor/block_buffer_36_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_35_s0  (
	.D(\top/processor/n11293_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [35])
);
defparam \top/processor/block_buffer_35_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_34_s0  (
	.D(\top/processor/n11294_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [34])
);
defparam \top/processor/block_buffer_34_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_33_s0  (
	.D(\top/processor/n11295_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [33])
);
defparam \top/processor/block_buffer_33_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_32_s0  (
	.D(\top/processor/n11296_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_39_8 ),
	.Q(\top/processor/block_buffer [32])
);
defparam \top/processor/block_buffer_32_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_31_s0  (
	.D(\top/processor/n11297_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [31])
);
defparam \top/processor/block_buffer_31_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_30_s0  (
	.D(\top/processor/n11298_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [30])
);
defparam \top/processor/block_buffer_30_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_29_s0  (
	.D(\top/processor/n11299_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [29])
);
defparam \top/processor/block_buffer_29_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_28_s0  (
	.D(\top/processor/n11300_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [28])
);
defparam \top/processor/block_buffer_28_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_27_s0  (
	.D(\top/processor/n11301_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [27])
);
defparam \top/processor/block_buffer_27_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_26_s0  (
	.D(\top/processor/n11302_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [26])
);
defparam \top/processor/block_buffer_26_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_25_s0  (
	.D(\top/processor/n11303_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [25])
);
defparam \top/processor/block_buffer_25_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_24_s0  (
	.D(\top/processor/n11304_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_31_8 ),
	.Q(\top/processor/block_buffer [24])
);
defparam \top/processor/block_buffer_24_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_23_s0  (
	.D(\top/processor/n11305_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [23])
);
defparam \top/processor/block_buffer_23_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_22_s0  (
	.D(\top/processor/n11306_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [22])
);
defparam \top/processor/block_buffer_22_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_21_s0  (
	.D(\top/processor/n11307_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [21])
);
defparam \top/processor/block_buffer_21_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_20_s0  (
	.D(\top/processor/n11308_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [20])
);
defparam \top/processor/block_buffer_20_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_19_s0  (
	.D(\top/processor/n11309_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [19])
);
defparam \top/processor/block_buffer_19_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_18_s0  (
	.D(\top/processor/n11310_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [18])
);
defparam \top/processor/block_buffer_18_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_17_s0  (
	.D(\top/processor/n11311_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [17])
);
defparam \top/processor/block_buffer_17_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_16_s0  (
	.D(\top/processor/n11312_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_23_8 ),
	.Q(\top/processor/block_buffer [16])
);
defparam \top/processor/block_buffer_16_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_15_s0  (
	.D(\top/processor/n11313_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [15])
);
defparam \top/processor/block_buffer_15_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_14_s0  (
	.D(\top/processor/n11314_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [14])
);
defparam \top/processor/block_buffer_14_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_13_s0  (
	.D(\top/processor/n11315_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [13])
);
defparam \top/processor/block_buffer_13_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_12_s0  (
	.D(\top/processor/n11316_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [12])
);
defparam \top/processor/block_buffer_12_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_11_s0  (
	.D(\top/processor/n11317_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [11])
);
defparam \top/processor/block_buffer_11_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_10_s0  (
	.D(\top/processor/n11318_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [10])
);
defparam \top/processor/block_buffer_10_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_9_s0  (
	.D(\top/processor/n11319_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [9])
);
defparam \top/processor/block_buffer_9_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_8_s0  (
	.D(\top/processor/n11320_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_15_8 ),
	.Q(\top/processor/block_buffer [8])
);
defparam \top/processor/block_buffer_8_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_7_s0  (
	.D(\top/processor/n11321_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [7])
);
defparam \top/processor/block_buffer_7_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_6_s0  (
	.D(\top/processor/n11322_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [6])
);
defparam \top/processor/block_buffer_6_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_5_s0  (
	.D(\top/processor/n11323_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [5])
);
defparam \top/processor/block_buffer_5_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_4_s0  (
	.D(\top/processor/n11324_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [4])
);
defparam \top/processor/block_buffer_4_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_3_s0  (
	.D(\top/processor/n11325_12 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [3])
);
defparam \top/processor/block_buffer_3_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_2_s0  (
	.D(\top/processor/n10822_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [2])
);
defparam \top/processor/block_buffer_2_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_1_s0  (
	.D(\top/processor/n10823_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [1])
);
defparam \top/processor/block_buffer_1_s0 .INIT=1'b0;
DFFE \top/processor/block_buffer_0_s0  (
	.D(\top/processor/n10824_15 ),
	.CLK(clk),
	.CE(\top/processor/block_buffer_7_11 ),
	.Q(\top/processor/block_buffer [0])
);
defparam \top/processor/block_buffer_0_s0 .INIT=1'b0;
DFFC \top/processor/state_2_s0  (
	.D(\top/processor/n11362_17 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/state_0 [2])
);
defparam \top/processor/state_2_s0 .INIT=1'b0;
DFFPE \top/processor/hash_state_254_s0  (
	.D(\top/processor/n10562_16 ),
	.CLK(clk),
	.CE(\top/processor/hash_state_255_7 ),
	.PRESET(rst),
	.Q(\top/hash_out [254])
);
defparam \top/processor/hash_state_254_s0 .INIT=1'b1;
DFFCE \top/processor/core_start_s1  (
	.D(\top/processor/n9789_16 ),
	.CLK(clk),
	.CE(\top/processor/core_start_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_start )
);
defparam \top/processor/core_start_s1 .INIT=1'b0;
LUT4 \top/processor/sha_core/n3494_s182  (
	.I0(\top/processor/sha_core/n3494_149 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_150 ),
	.I3(\top/processor/sha_core/n3494_151 ),
	.F(\top/processor/sha_core/n3494_148 )
);
defparam \top/processor/sha_core/n3494_s182 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3866_s134  (
	.I0(\top/processor/sha_core/n3866_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_117 ),
	.I3(\top/processor/sha_core/n3494_151 ),
	.F(\top/processor/sha_core/n3866_101 )
);
defparam \top/processor/sha_core/n3866_s134 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3705_s143  (
	.I0(\top/processor/sha_core/n3607_164 ),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[34] [31]),
	.I3(\top/processor/sha_core/w[35] [31]),
	.F(\top/processor/sha_core/n3607_133 )
);
defparam \top/processor/sha_core/n3705_s143 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3706_s143  (
	.I0(\top/processor/sha_core/n3608_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [30]),
	.I3(\top/processor/sha_core/w[32] [30]),
	.F(\top/processor/sha_core/n3608_133 )
);
defparam \top/processor/sha_core/n3706_s143 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3707_s143  (
	.I0(\top/processor/sha_core/n3609_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [29]),
	.I3(\top/processor/sha_core/w[32] [29]),
	.F(\top/processor/sha_core/n3609_133 )
);
defparam \top/processor/sha_core/n3707_s143 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3708_s143  (
	.I0(\top/processor/sha_core/n3610_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [28]),
	.I3(\top/processor/sha_core/w[32] [28]),
	.F(\top/processor/sha_core/n3610_133 )
);
defparam \top/processor/sha_core/n3708_s143 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3709_s143  (
	.I0(\top/processor/sha_core/n3611_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [27]),
	.I3(\top/processor/sha_core/w[32] [27]),
	.F(\top/processor/sha_core/n3611_133 )
);
defparam \top/processor/sha_core/n3709_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s143  (
	.I0(\top/processor/sha_core/n3612_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [26]),
	.I3(\top/processor/sha_core/w[32] [26]),
	.F(\top/processor/sha_core/n3612_133 )
);
defparam \top/processor/sha_core/n3710_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s143  (
	.I0(\top/processor/sha_core/n3613_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [25]),
	.I3(\top/processor/sha_core/w[32] [25]),
	.F(\top/processor/sha_core/n3613_133 )
);
defparam \top/processor/sha_core/n3711_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s143  (
	.I0(\top/processor/sha_core/n3614_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [24]),
	.I3(\top/processor/sha_core/w[32] [24]),
	.F(\top/processor/sha_core/n3614_133 )
);
defparam \top/processor/sha_core/n3712_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s143  (
	.I0(\top/processor/sha_core/n3615_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [23]),
	.I3(\top/processor/sha_core/w[32] [23]),
	.F(\top/processor/sha_core/n3615_133 )
);
defparam \top/processor/sha_core/n3713_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s143  (
	.I0(\top/processor/sha_core/n3616_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [22]),
	.I3(\top/processor/sha_core/w[32] [22]),
	.F(\top/processor/sha_core/n3616_133 )
);
defparam \top/processor/sha_core/n3714_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s143  (
	.I0(\top/processor/sha_core/n3617_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [21]),
	.I3(\top/processor/sha_core/w[32] [21]),
	.F(\top/processor/sha_core/n3617_133 )
);
defparam \top/processor/sha_core/n3715_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s143  (
	.I0(\top/processor/sha_core/n3618_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [20]),
	.I3(\top/processor/sha_core/w[32] [20]),
	.F(\top/processor/sha_core/n3618_133 )
);
defparam \top/processor/sha_core/n3716_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s143  (
	.I0(\top/processor/sha_core/n3619_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [19]),
	.I3(\top/processor/sha_core/w[32] [19]),
	.F(\top/processor/sha_core/n3619_133 )
);
defparam \top/processor/sha_core/n3717_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s143  (
	.I0(\top/processor/sha_core/n3620_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [18]),
	.I3(\top/processor/sha_core/w[32] [18]),
	.F(\top/processor/sha_core/n3620_133 )
);
defparam \top/processor/sha_core/n3718_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s143  (
	.I0(\top/processor/sha_core/n3621_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [17]),
	.I3(\top/processor/sha_core/w[32] [17]),
	.F(\top/processor/sha_core/n3621_133 )
);
defparam \top/processor/sha_core/n3719_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s183  (
	.I0(\top/processor/sha_core/n3494_152 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_153 ),
	.I3(\top/processor/sha_core/n3494_154 ),
	.F(\top/processor/sha_core/n3494_135 )
);
defparam \top/processor/sha_core/n3494_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s135  (
	.I0(\top/processor/sha_core/n3866_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_119 ),
	.I3(\top/processor/sha_core/n3494_154 ),
	.F(\top/processor/sha_core/n3866_103 )
);
defparam \top/processor/sha_core/n3866_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3720_s143  (
	.I0(\top/processor/sha_core/n3622_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [16]),
	.I3(\top/processor/sha_core/w[32] [16]),
	.F(\top/processor/sha_core/n3622_133 )
);
defparam \top/processor/sha_core/n3720_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s143  (
	.I0(\top/processor/sha_core/n3623_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [15]),
	.I3(\top/processor/sha_core/w[32] [15]),
	.F(\top/processor/sha_core/n3623_133 )
);
defparam \top/processor/sha_core/n3721_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s143  (
	.I0(\top/processor/sha_core/n3624_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [14]),
	.I3(\top/processor/sha_core/w[32] [14]),
	.F(\top/processor/sha_core/n3624_133 )
);
defparam \top/processor/sha_core/n3722_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s143  (
	.I0(\top/processor/sha_core/n3625_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [13]),
	.I3(\top/processor/sha_core/w[32] [13]),
	.F(\top/processor/sha_core/n3625_133 )
);
defparam \top/processor/sha_core/n3723_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s143  (
	.I0(\top/processor/sha_core/n3626_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [12]),
	.I3(\top/processor/sha_core/w[32] [12]),
	.F(\top/processor/sha_core/n3626_133 )
);
defparam \top/processor/sha_core/n3724_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s143  (
	.I0(\top/processor/sha_core/n3627_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [11]),
	.I3(\top/processor/sha_core/w[32] [11]),
	.F(\top/processor/sha_core/n3627_133 )
);
defparam \top/processor/sha_core/n3725_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s143  (
	.I0(\top/processor/sha_core/n3628_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [10]),
	.I3(\top/processor/sha_core/w[32] [10]),
	.F(\top/processor/sha_core/n3628_133 )
);
defparam \top/processor/sha_core/n3726_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s143  (
	.I0(\top/processor/sha_core/n3629_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [9]),
	.I3(\top/processor/sha_core/w[32] [9]),
	.F(\top/processor/sha_core/n3629_133 )
);
defparam \top/processor/sha_core/n3727_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s143  (
	.I0(\top/processor/sha_core/n3630_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [8]),
	.I3(\top/processor/sha_core/w[32] [8]),
	.F(\top/processor/sha_core/n3630_133 )
);
defparam \top/processor/sha_core/n3728_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s143  (
	.I0(\top/processor/sha_core/n3631_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [7]),
	.I3(\top/processor/sha_core/w[32] [7]),
	.F(\top/processor/sha_core/n3631_133 )
);
defparam \top/processor/sha_core/n3729_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s143  (
	.I0(\top/processor/sha_core/n3632_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [6]),
	.I3(\top/processor/sha_core/w[32] [6]),
	.F(\top/processor/sha_core/n3632_133 )
);
defparam \top/processor/sha_core/n3730_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s143  (
	.I0(\top/processor/sha_core/n3633_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [5]),
	.I3(\top/processor/sha_core/w[32] [5]),
	.F(\top/processor/sha_core/n3633_133 )
);
defparam \top/processor/sha_core/n3731_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s143  (
	.I0(\top/processor/sha_core/n3634_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [4]),
	.I3(\top/processor/sha_core/w[32] [4]),
	.F(\top/processor/sha_core/n3634_133 )
);
defparam \top/processor/sha_core/n3732_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s143  (
	.I0(\top/processor/sha_core/n3635_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [3]),
	.I3(\top/processor/sha_core/w[32] [3]),
	.F(\top/processor/sha_core/n3635_133 )
);
defparam \top/processor/sha_core/n3733_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s143  (
	.I0(\top/processor/sha_core/n3636_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [2]),
	.I3(\top/processor/sha_core/w[32] [2]),
	.F(\top/processor/sha_core/n3636_133 )
);
defparam \top/processor/sha_core/n3734_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s143  (
	.I0(\top/processor/sha_core/n3637_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [1]),
	.I3(\top/processor/sha_core/w[32] [1]),
	.F(\top/processor/sha_core/n3637_133 )
);
defparam \top/processor/sha_core/n3735_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s143  (
	.I0(\top/processor/sha_core/n3638_164 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[34] [0]),
	.I3(\top/processor/sha_core/w[32] [0]),
	.F(\top/processor/sha_core/n3638_133 )
);
defparam \top/processor/sha_core/n3736_s143 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s184  (
	.I0(\top/processor/sha_core/n3494_155 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_156 ),
	.I3(\top/processor/sha_core/n3494_157 ),
	.F(\top/processor/sha_core/n3494_137 )
);
defparam \top/processor/sha_core/n3494_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s136  (
	.I0(\top/processor/sha_core/n3866_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_121 ),
	.I3(\top/processor/sha_core/n3494_157 ),
	.F(\top/processor/sha_core/n3866_105 )
);
defparam \top/processor/sha_core/n3866_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3494_s185  (
	.I0(\top/processor/sha_core/n3494_158 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_159 ),
	.I3(\top/processor/sha_core/n3494_160 ),
	.F(\top/processor/sha_core/n3494_139 )
);
defparam \top/processor/sha_core/n3494_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s137  (
	.I0(\top/processor/sha_core/n3866_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_123 ),
	.I3(\top/processor/sha_core/n3494_160 ),
	.F(\top/processor/sha_core/n3866_107 )
);
defparam \top/processor/sha_core/n3866_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s144  (
	.I0(\top/processor/sha_core/n3607_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [31]),
	.I3(\top/processor/sha_core/w[36] [31]),
	.F(\top/processor/sha_core/n3607_135 )
);
defparam \top/processor/sha_core/n3705_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s144  (
	.I0(\top/processor/sha_core/n3608_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [30]),
	.I3(\top/processor/sha_core/w[36] [30]),
	.F(\top/processor/sha_core/n3608_135 )
);
defparam \top/processor/sha_core/n3706_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s144  (
	.I0(\top/processor/sha_core/n3609_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [29]),
	.I3(\top/processor/sha_core/w[36] [29]),
	.F(\top/processor/sha_core/n3609_135 )
);
defparam \top/processor/sha_core/n3707_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s144  (
	.I0(\top/processor/sha_core/n3610_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [28]),
	.I3(\top/processor/sha_core/w[36] [28]),
	.F(\top/processor/sha_core/n3610_135 )
);
defparam \top/processor/sha_core/n3708_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s144  (
	.I0(\top/processor/sha_core/n3611_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [27]),
	.I3(\top/processor/sha_core/w[36] [27]),
	.F(\top/processor/sha_core/n3611_135 )
);
defparam \top/processor/sha_core/n3709_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s144  (
	.I0(\top/processor/sha_core/n3612_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [26]),
	.I3(\top/processor/sha_core/w[36] [26]),
	.F(\top/processor/sha_core/n3612_135 )
);
defparam \top/processor/sha_core/n3710_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s144  (
	.I0(\top/processor/sha_core/n3613_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [25]),
	.I3(\top/processor/sha_core/w[36] [25]),
	.F(\top/processor/sha_core/n3613_135 )
);
defparam \top/processor/sha_core/n3711_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s144  (
	.I0(\top/processor/sha_core/n3614_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [24]),
	.I3(\top/processor/sha_core/w[36] [24]),
	.F(\top/processor/sha_core/n3614_135 )
);
defparam \top/processor/sha_core/n3712_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s144  (
	.I0(\top/processor/sha_core/n3615_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [23]),
	.I3(\top/processor/sha_core/w[36] [23]),
	.F(\top/processor/sha_core/n3615_135 )
);
defparam \top/processor/sha_core/n3713_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s144  (
	.I0(\top/processor/sha_core/n3616_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [22]),
	.I3(\top/processor/sha_core/w[36] [22]),
	.F(\top/processor/sha_core/n3616_135 )
);
defparam \top/processor/sha_core/n3714_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s144  (
	.I0(\top/processor/sha_core/n3617_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [21]),
	.I3(\top/processor/sha_core/w[36] [21]),
	.F(\top/processor/sha_core/n3617_135 )
);
defparam \top/processor/sha_core/n3715_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s186  (
	.I0(\top/processor/sha_core/n3494_161 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_162 ),
	.I3(\top/processor/sha_core/n3494_163 ),
	.F(\top/processor/sha_core/n3494_141 )
);
defparam \top/processor/sha_core/n3494_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s138  (
	.I0(\top/processor/sha_core/n3866_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_125 ),
	.I3(\top/processor/sha_core/n3494_163 ),
	.F(\top/processor/sha_core/n3866_109 )
);
defparam \top/processor/sha_core/n3866_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3716_s144  (
	.I0(\top/processor/sha_core/n3618_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [20]),
	.I3(\top/processor/sha_core/w[36] [20]),
	.F(\top/processor/sha_core/n3618_135 )
);
defparam \top/processor/sha_core/n3716_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s144  (
	.I0(\top/processor/sha_core/n3619_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [19]),
	.I3(\top/processor/sha_core/w[36] [19]),
	.F(\top/processor/sha_core/n3619_135 )
);
defparam \top/processor/sha_core/n3717_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s144  (
	.I0(\top/processor/sha_core/n3620_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [18]),
	.I3(\top/processor/sha_core/w[36] [18]),
	.F(\top/processor/sha_core/n3620_135 )
);
defparam \top/processor/sha_core/n3718_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s144  (
	.I0(\top/processor/sha_core/n3621_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [17]),
	.I3(\top/processor/sha_core/w[36] [17]),
	.F(\top/processor/sha_core/n3621_135 )
);
defparam \top/processor/sha_core/n3719_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s144  (
	.I0(\top/processor/sha_core/n3622_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [16]),
	.I3(\top/processor/sha_core/w[36] [16]),
	.F(\top/processor/sha_core/n3622_135 )
);
defparam \top/processor/sha_core/n3720_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s144  (
	.I0(\top/processor/sha_core/n3623_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [15]),
	.I3(\top/processor/sha_core/w[36] [15]),
	.F(\top/processor/sha_core/n3623_135 )
);
defparam \top/processor/sha_core/n3721_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s144  (
	.I0(\top/processor/sha_core/n3624_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [14]),
	.I3(\top/processor/sha_core/w[36] [14]),
	.F(\top/processor/sha_core/n3624_135 )
);
defparam \top/processor/sha_core/n3722_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s144  (
	.I0(\top/processor/sha_core/n3625_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [13]),
	.I3(\top/processor/sha_core/w[36] [13]),
	.F(\top/processor/sha_core/n3625_135 )
);
defparam \top/processor/sha_core/n3723_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s144  (
	.I0(\top/processor/sha_core/n3626_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [12]),
	.I3(\top/processor/sha_core/w[36] [12]),
	.F(\top/processor/sha_core/n3626_135 )
);
defparam \top/processor/sha_core/n3724_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s144  (
	.I0(\top/processor/sha_core/n3627_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [11]),
	.I3(\top/processor/sha_core/w[36] [11]),
	.F(\top/processor/sha_core/n3627_135 )
);
defparam \top/processor/sha_core/n3725_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s144  (
	.I0(\top/processor/sha_core/n3628_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [10]),
	.I3(\top/processor/sha_core/w[36] [10]),
	.F(\top/processor/sha_core/n3628_135 )
);
defparam \top/processor/sha_core/n3726_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s144  (
	.I0(\top/processor/sha_core/n3629_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [9]),
	.I3(\top/processor/sha_core/w[36] [9]),
	.F(\top/processor/sha_core/n3629_135 )
);
defparam \top/processor/sha_core/n3727_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s144  (
	.I0(\top/processor/sha_core/n3630_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [8]),
	.I3(\top/processor/sha_core/w[36] [8]),
	.F(\top/processor/sha_core/n3630_135 )
);
defparam \top/processor/sha_core/n3728_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s144  (
	.I0(\top/processor/sha_core/n3631_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [7]),
	.I3(\top/processor/sha_core/w[36] [7]),
	.F(\top/processor/sha_core/n3631_135 )
);
defparam \top/processor/sha_core/n3729_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s144  (
	.I0(\top/processor/sha_core/n3632_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [6]),
	.I3(\top/processor/sha_core/w[36] [6]),
	.F(\top/processor/sha_core/n3632_135 )
);
defparam \top/processor/sha_core/n3730_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s144  (
	.I0(\top/processor/sha_core/n3633_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [5]),
	.I3(\top/processor/sha_core/w[36] [5]),
	.F(\top/processor/sha_core/n3633_135 )
);
defparam \top/processor/sha_core/n3731_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s144  (
	.I0(\top/processor/sha_core/n3634_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [4]),
	.I3(\top/processor/sha_core/w[36] [4]),
	.F(\top/processor/sha_core/n3634_135 )
);
defparam \top/processor/sha_core/n3732_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s144  (
	.I0(\top/processor/sha_core/n3635_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [3]),
	.I3(\top/processor/sha_core/w[36] [3]),
	.F(\top/processor/sha_core/n3635_135 )
);
defparam \top/processor/sha_core/n3733_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s144  (
	.I0(\top/processor/sha_core/n3636_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [2]),
	.I3(\top/processor/sha_core/w[36] [2]),
	.F(\top/processor/sha_core/n3636_135 )
);
defparam \top/processor/sha_core/n3734_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s144  (
	.I0(\top/processor/sha_core/n3637_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [1]),
	.I3(\top/processor/sha_core/w[36] [1]),
	.F(\top/processor/sha_core/n3637_135 )
);
defparam \top/processor/sha_core/n3735_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s187  (
	.I0(\top/processor/sha_core/n3494_164 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_165 ),
	.I3(\top/processor/sha_core/n3494_166 ),
	.F(\top/processor/sha_core/n3494_143 )
);
defparam \top/processor/sha_core/n3494_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s139  (
	.I0(\top/processor/sha_core/n3866_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_127 ),
	.I3(\top/processor/sha_core/n3494_166 ),
	.F(\top/processor/sha_core/n3866_111 )
);
defparam \top/processor/sha_core/n3866_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3736_s144  (
	.I0(\top/processor/sha_core/n3638_165 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[38] [0]),
	.I3(\top/processor/sha_core/w[36] [0]),
	.F(\top/processor/sha_core/n3638_135 )
);
defparam \top/processor/sha_core/n3736_s144 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s180  (
	.I0(\top/processor/sha_core/n3495_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_149 ),
	.I3(\top/processor/sha_core/n3495_150 ),
	.F(\top/processor/sha_core/n3495_133 )
);
defparam \top/processor/sha_core/n3495_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s132  (
	.I0(\top/processor/sha_core/n3867_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_117 ),
	.I3(\top/processor/sha_core/n3495_150 ),
	.F(\top/processor/sha_core/n3867_101 )
);
defparam \top/processor/sha_core/n3867_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s145  (
	.I0(\top/processor/sha_core/n3607_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [31]),
	.I3(\top/processor/sha_core/w[40] [31]),
	.F(\top/processor/sha_core/n3607_137 )
);
defparam \top/processor/sha_core/n3705_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s145  (
	.I0(\top/processor/sha_core/n3608_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [30]),
	.I3(\top/processor/sha_core/w[40] [30]),
	.F(\top/processor/sha_core/n3608_137 )
);
defparam \top/processor/sha_core/n3706_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s145  (
	.I0(\top/processor/sha_core/n3609_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [29]),
	.I3(\top/processor/sha_core/w[40] [29]),
	.F(\top/processor/sha_core/n3609_137 )
);
defparam \top/processor/sha_core/n3707_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s145  (
	.I0(\top/processor/sha_core/n3610_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [28]),
	.I3(\top/processor/sha_core/w[40] [28]),
	.F(\top/processor/sha_core/n3610_137 )
);
defparam \top/processor/sha_core/n3708_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s145  (
	.I0(\top/processor/sha_core/n3611_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [27]),
	.I3(\top/processor/sha_core/w[40] [27]),
	.F(\top/processor/sha_core/n3611_137 )
);
defparam \top/processor/sha_core/n3709_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s145  (
	.I0(\top/processor/sha_core/n3612_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [26]),
	.I3(\top/processor/sha_core/w[40] [26]),
	.F(\top/processor/sha_core/n3612_137 )
);
defparam \top/processor/sha_core/n3710_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s145  (
	.I0(\top/processor/sha_core/n3613_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [25]),
	.I3(\top/processor/sha_core/w[40] [25]),
	.F(\top/processor/sha_core/n3613_137 )
);
defparam \top/processor/sha_core/n3711_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s181  (
	.I0(\top/processor/sha_core/n3495_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_152 ),
	.I3(\top/processor/sha_core/n3495_153 ),
	.F(\top/processor/sha_core/n3495_135 )
);
defparam \top/processor/sha_core/n3495_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s133  (
	.I0(\top/processor/sha_core/n3867_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_119 ),
	.I3(\top/processor/sha_core/n3495_153 ),
	.F(\top/processor/sha_core/n3867_103 )
);
defparam \top/processor/sha_core/n3867_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3712_s145  (
	.I0(\top/processor/sha_core/n3614_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [24]),
	.I3(\top/processor/sha_core/w[40] [24]),
	.F(\top/processor/sha_core/n3614_137 )
);
defparam \top/processor/sha_core/n3712_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s145  (
	.I0(\top/processor/sha_core/n3615_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [23]),
	.I3(\top/processor/sha_core/w[40] [23]),
	.F(\top/processor/sha_core/n3615_137 )
);
defparam \top/processor/sha_core/n3713_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s145  (
	.I0(\top/processor/sha_core/n3616_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [22]),
	.I3(\top/processor/sha_core/w[40] [22]),
	.F(\top/processor/sha_core/n3616_137 )
);
defparam \top/processor/sha_core/n3714_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s145  (
	.I0(\top/processor/sha_core/n3617_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [21]),
	.I3(\top/processor/sha_core/w[40] [21]),
	.F(\top/processor/sha_core/n3617_137 )
);
defparam \top/processor/sha_core/n3715_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s145  (
	.I0(\top/processor/sha_core/n3618_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [20]),
	.I3(\top/processor/sha_core/w[40] [20]),
	.F(\top/processor/sha_core/n3618_137 )
);
defparam \top/processor/sha_core/n3716_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s145  (
	.I0(\top/processor/sha_core/n3619_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [19]),
	.I3(\top/processor/sha_core/w[40] [19]),
	.F(\top/processor/sha_core/n3619_137 )
);
defparam \top/processor/sha_core/n3717_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s145  (
	.I0(\top/processor/sha_core/n3620_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [18]),
	.I3(\top/processor/sha_core/w[40] [18]),
	.F(\top/processor/sha_core/n3620_137 )
);
defparam \top/processor/sha_core/n3718_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s145  (
	.I0(\top/processor/sha_core/n3621_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [17]),
	.I3(\top/processor/sha_core/w[40] [17]),
	.F(\top/processor/sha_core/n3621_137 )
);
defparam \top/processor/sha_core/n3719_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s145  (
	.I0(\top/processor/sha_core/n3622_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [16]),
	.I3(\top/processor/sha_core/w[40] [16]),
	.F(\top/processor/sha_core/n3622_137 )
);
defparam \top/processor/sha_core/n3720_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s145  (
	.I0(\top/processor/sha_core/n3623_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [15]),
	.I3(\top/processor/sha_core/w[40] [15]),
	.F(\top/processor/sha_core/n3623_137 )
);
defparam \top/processor/sha_core/n3721_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s145  (
	.I0(\top/processor/sha_core/n3624_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [14]),
	.I3(\top/processor/sha_core/w[40] [14]),
	.F(\top/processor/sha_core/n3624_137 )
);
defparam \top/processor/sha_core/n3722_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s145  (
	.I0(\top/processor/sha_core/n3625_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [13]),
	.I3(\top/processor/sha_core/w[40] [13]),
	.F(\top/processor/sha_core/n3625_137 )
);
defparam \top/processor/sha_core/n3723_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s145  (
	.I0(\top/processor/sha_core/n3626_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [12]),
	.I3(\top/processor/sha_core/w[40] [12]),
	.F(\top/processor/sha_core/n3626_137 )
);
defparam \top/processor/sha_core/n3724_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s145  (
	.I0(\top/processor/sha_core/n3627_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [11]),
	.I3(\top/processor/sha_core/w[40] [11]),
	.F(\top/processor/sha_core/n3627_137 )
);
defparam \top/processor/sha_core/n3725_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s145  (
	.I0(\top/processor/sha_core/n3628_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [10]),
	.I3(\top/processor/sha_core/w[40] [10]),
	.F(\top/processor/sha_core/n3628_137 )
);
defparam \top/processor/sha_core/n3726_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s145  (
	.I0(\top/processor/sha_core/n3629_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [9]),
	.I3(\top/processor/sha_core/w[40] [9]),
	.F(\top/processor/sha_core/n3629_137 )
);
defparam \top/processor/sha_core/n3727_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s145  (
	.I0(\top/processor/sha_core/n3630_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [8]),
	.I3(\top/processor/sha_core/w[40] [8]),
	.F(\top/processor/sha_core/n3630_137 )
);
defparam \top/processor/sha_core/n3728_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s145  (
	.I0(\top/processor/sha_core/n3631_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [7]),
	.I3(\top/processor/sha_core/w[40] [7]),
	.F(\top/processor/sha_core/n3631_137 )
);
defparam \top/processor/sha_core/n3729_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s145  (
	.I0(\top/processor/sha_core/n3632_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [6]),
	.I3(\top/processor/sha_core/w[40] [6]),
	.F(\top/processor/sha_core/n3632_137 )
);
defparam \top/processor/sha_core/n3730_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s145  (
	.I0(\top/processor/sha_core/n3633_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [5]),
	.I3(\top/processor/sha_core/w[40] [5]),
	.F(\top/processor/sha_core/n3633_137 )
);
defparam \top/processor/sha_core/n3731_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s182  (
	.I0(\top/processor/sha_core/n3495_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_155 ),
	.I3(\top/processor/sha_core/n3495_156 ),
	.F(\top/processor/sha_core/n3495_137 )
);
defparam \top/processor/sha_core/n3495_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s134  (
	.I0(\top/processor/sha_core/n3867_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_121 ),
	.I3(\top/processor/sha_core/n3495_156 ),
	.F(\top/processor/sha_core/n3867_105 )
);
defparam \top/processor/sha_core/n3867_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3732_s145  (
	.I0(\top/processor/sha_core/n3634_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [4]),
	.I3(\top/processor/sha_core/w[40] [4]),
	.F(\top/processor/sha_core/n3634_137 )
);
defparam \top/processor/sha_core/n3732_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s145  (
	.I0(\top/processor/sha_core/n3635_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [3]),
	.I3(\top/processor/sha_core/w[40] [3]),
	.F(\top/processor/sha_core/n3635_137 )
);
defparam \top/processor/sha_core/n3733_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s145  (
	.I0(\top/processor/sha_core/n3636_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [2]),
	.I3(\top/processor/sha_core/w[40] [2]),
	.F(\top/processor/sha_core/n3636_137 )
);
defparam \top/processor/sha_core/n3734_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s145  (
	.I0(\top/processor/sha_core/n3637_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [1]),
	.I3(\top/processor/sha_core/w[40] [1]),
	.F(\top/processor/sha_core/n3637_137 )
);
defparam \top/processor/sha_core/n3735_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s145  (
	.I0(\top/processor/sha_core/n3638_166 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[42] [0]),
	.I3(\top/processor/sha_core/w[40] [0]),
	.F(\top/processor/sha_core/n3638_137 )
);
defparam \top/processor/sha_core/n3736_s145 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s183  (
	.I0(\top/processor/sha_core/n3495_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_158 ),
	.I3(\top/processor/sha_core/n3495_159 ),
	.F(\top/processor/sha_core/n3495_139 )
);
defparam \top/processor/sha_core/n3495_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s135  (
	.I0(\top/processor/sha_core/n3867_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_123 ),
	.I3(\top/processor/sha_core/n3495_159 ),
	.F(\top/processor/sha_core/n3867_107 )
);
defparam \top/processor/sha_core/n3867_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s185  (
	.I0(\top/processor/sha_core/n3488_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_149 ),
	.I3(\top/processor/sha_core/n3488_150 ),
	.F(\top/processor/sha_core/n3488_133 )
);
defparam \top/processor/sha_core/n3488_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s137  (
	.I0(\top/processor/sha_core/n3860_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_117 ),
	.I3(\top/processor/sha_core/n3488_150 ),
	.F(\top/processor/sha_core/n3860_101 )
);
defparam \top/processor/sha_core/n3860_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s146  (
	.I0(\top/processor/sha_core/n3607_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [31]),
	.I3(\top/processor/sha_core/w[44] [31]),
	.F(\top/processor/sha_core/n3607_139 )
);
defparam \top/processor/sha_core/n3705_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s146  (
	.I0(\top/processor/sha_core/n3608_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [30]),
	.I3(\top/processor/sha_core/w[44] [30]),
	.F(\top/processor/sha_core/n3608_139 )
);
defparam \top/processor/sha_core/n3706_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s146  (
	.I0(\top/processor/sha_core/n3609_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [29]),
	.I3(\top/processor/sha_core/w[44] [29]),
	.F(\top/processor/sha_core/n3609_139 )
);
defparam \top/processor/sha_core/n3707_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s184  (
	.I0(\top/processor/sha_core/n3495_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_161 ),
	.I3(\top/processor/sha_core/n3495_162 ),
	.F(\top/processor/sha_core/n3495_141 )
);
defparam \top/processor/sha_core/n3495_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s136  (
	.I0(\top/processor/sha_core/n3867_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_125 ),
	.I3(\top/processor/sha_core/n3495_162 ),
	.F(\top/processor/sha_core/n3867_109 )
);
defparam \top/processor/sha_core/n3867_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3708_s146  (
	.I0(\top/processor/sha_core/n3610_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [28]),
	.I3(\top/processor/sha_core/w[44] [28]),
	.F(\top/processor/sha_core/n3610_139 )
);
defparam \top/processor/sha_core/n3708_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s146  (
	.I0(\top/processor/sha_core/n3611_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [27]),
	.I3(\top/processor/sha_core/w[44] [27]),
	.F(\top/processor/sha_core/n3611_139 )
);
defparam \top/processor/sha_core/n3709_s146 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3710_s146  (
	.I0(\top/processor/sha_core/n3612_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [26]),
	.I3(\top/processor/sha_core/w[44] [26]),
	.F(\top/processor/sha_core/n3612_139 )
);
defparam \top/processor/sha_core/n3710_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s146  (
	.I0(\top/processor/sha_core/n3613_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [25]),
	.I3(\top/processor/sha_core/w[44] [25]),
	.F(\top/processor/sha_core/n3613_139 )
);
defparam \top/processor/sha_core/n3711_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s146  (
	.I0(\top/processor/sha_core/n3614_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [24]),
	.I3(\top/processor/sha_core/w[44] [24]),
	.F(\top/processor/sha_core/n3614_139 )
);
defparam \top/processor/sha_core/n3712_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s146  (
	.I0(\top/processor/sha_core/n3615_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [23]),
	.I3(\top/processor/sha_core/w[44] [23]),
	.F(\top/processor/sha_core/n3615_139 )
);
defparam \top/processor/sha_core/n3713_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s146  (
	.I0(\top/processor/sha_core/n3616_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [22]),
	.I3(\top/processor/sha_core/w[44] [22]),
	.F(\top/processor/sha_core/n3616_139 )
);
defparam \top/processor/sha_core/n3714_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s146  (
	.I0(\top/processor/sha_core/n3617_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [21]),
	.I3(\top/processor/sha_core/w[44] [21]),
	.F(\top/processor/sha_core/n3617_139 )
);
defparam \top/processor/sha_core/n3715_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s146  (
	.I0(\top/processor/sha_core/n3618_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [20]),
	.I3(\top/processor/sha_core/w[44] [20]),
	.F(\top/processor/sha_core/n3618_139 )
);
defparam \top/processor/sha_core/n3716_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s146  (
	.I0(\top/processor/sha_core/n3619_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [19]),
	.I3(\top/processor/sha_core/w[44] [19]),
	.F(\top/processor/sha_core/n3619_139 )
);
defparam \top/processor/sha_core/n3717_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s146  (
	.I0(\top/processor/sha_core/n3620_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [18]),
	.I3(\top/processor/sha_core/w[44] [18]),
	.F(\top/processor/sha_core/n3620_139 )
);
defparam \top/processor/sha_core/n3718_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s146  (
	.I0(\top/processor/sha_core/n3621_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [17]),
	.I3(\top/processor/sha_core/w[44] [17]),
	.F(\top/processor/sha_core/n3621_139 )
);
defparam \top/processor/sha_core/n3719_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s146  (
	.I0(\top/processor/sha_core/n3622_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [16]),
	.I3(\top/processor/sha_core/w[44] [16]),
	.F(\top/processor/sha_core/n3622_139 )
);
defparam \top/processor/sha_core/n3720_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s146  (
	.I0(\top/processor/sha_core/n3623_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [15]),
	.I3(\top/processor/sha_core/w[44] [15]),
	.F(\top/processor/sha_core/n3623_139 )
);
defparam \top/processor/sha_core/n3721_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s146  (
	.I0(\top/processor/sha_core/n3624_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [14]),
	.I3(\top/processor/sha_core/w[44] [14]),
	.F(\top/processor/sha_core/n3624_139 )
);
defparam \top/processor/sha_core/n3722_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s146  (
	.I0(\top/processor/sha_core/n3625_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [13]),
	.I3(\top/processor/sha_core/w[44] [13]),
	.F(\top/processor/sha_core/n3625_139 )
);
defparam \top/processor/sha_core/n3723_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s146  (
	.I0(\top/processor/sha_core/n3626_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [12]),
	.I3(\top/processor/sha_core/w[44] [12]),
	.F(\top/processor/sha_core/n3626_139 )
);
defparam \top/processor/sha_core/n3724_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s146  (
	.I0(\top/processor/sha_core/n3627_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [11]),
	.I3(\top/processor/sha_core/w[44] [11]),
	.F(\top/processor/sha_core/n3627_139 )
);
defparam \top/processor/sha_core/n3725_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s146  (
	.I0(\top/processor/sha_core/n3628_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [10]),
	.I3(\top/processor/sha_core/w[44] [10]),
	.F(\top/processor/sha_core/n3628_139 )
);
defparam \top/processor/sha_core/n3726_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s146  (
	.I0(\top/processor/sha_core/n3629_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [9]),
	.I3(\top/processor/sha_core/w[44] [9]),
	.F(\top/processor/sha_core/n3629_139 )
);
defparam \top/processor/sha_core/n3727_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s185  (
	.I0(\top/processor/sha_core/n3495_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_164 ),
	.I3(\top/processor/sha_core/n3495_165 ),
	.F(\top/processor/sha_core/n3495_143 )
);
defparam \top/processor/sha_core/n3495_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s137  (
	.I0(\top/processor/sha_core/n3867_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_127 ),
	.I3(\top/processor/sha_core/n3495_165 ),
	.F(\top/processor/sha_core/n3867_111 )
);
defparam \top/processor/sha_core/n3867_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3728_s146  (
	.I0(\top/processor/sha_core/n3630_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [8]),
	.I3(\top/processor/sha_core/w[44] [8]),
	.F(\top/processor/sha_core/n3630_139 )
);
defparam \top/processor/sha_core/n3728_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s146  (
	.I0(\top/processor/sha_core/n3631_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [7]),
	.I3(\top/processor/sha_core/w[44] [7]),
	.F(\top/processor/sha_core/n3631_139 )
);
defparam \top/processor/sha_core/n3729_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s146  (
	.I0(\top/processor/sha_core/n3632_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [6]),
	.I3(\top/processor/sha_core/w[44] [6]),
	.F(\top/processor/sha_core/n3632_139 )
);
defparam \top/processor/sha_core/n3730_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s146  (
	.I0(\top/processor/sha_core/n3633_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [5]),
	.I3(\top/processor/sha_core/w[44] [5]),
	.F(\top/processor/sha_core/n3633_139 )
);
defparam \top/processor/sha_core/n3731_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s146  (
	.I0(\top/processor/sha_core/n3634_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [4]),
	.I3(\top/processor/sha_core/w[44] [4]),
	.F(\top/processor/sha_core/n3634_139 )
);
defparam \top/processor/sha_core/n3732_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s146  (
	.I0(\top/processor/sha_core/n3635_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [3]),
	.I3(\top/processor/sha_core/w[44] [3]),
	.F(\top/processor/sha_core/n3635_139 )
);
defparam \top/processor/sha_core/n3733_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s146  (
	.I0(\top/processor/sha_core/n3636_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [2]),
	.I3(\top/processor/sha_core/w[44] [2]),
	.F(\top/processor/sha_core/n3636_139 )
);
defparam \top/processor/sha_core/n3734_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s146  (
	.I0(\top/processor/sha_core/n3637_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [1]),
	.I3(\top/processor/sha_core/w[44] [1]),
	.F(\top/processor/sha_core/n3637_139 )
);
defparam \top/processor/sha_core/n3735_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s146  (
	.I0(\top/processor/sha_core/n3638_167 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[46] [0]),
	.I3(\top/processor/sha_core/w[44] [0]),
	.F(\top/processor/sha_core/n3638_139 )
);
defparam \top/processor/sha_core/n3736_s146 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3495_s186  (
	.I0(\top/processor/sha_core/n3495_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_167 ),
	.I3(\top/processor/sha_core/n3495_168 ),
	.F(\top/processor/sha_core/n3495_145 )
);
defparam \top/processor/sha_core/n3495_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s138  (
	.I0(\top/processor/sha_core/n3867_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_129 ),
	.I3(\top/processor/sha_core/n3495_168 ),
	.F(\top/processor/sha_core/n3867_113 )
);
defparam \top/processor/sha_core/n3867_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3495_s187  (
	.I0(\top/processor/sha_core/n3495_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_170 ),
	.I3(\top/processor/sha_core/n3495_171 ),
	.F(\top/processor/sha_core/n3495_147 )
);
defparam \top/processor/sha_core/n3495_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3867_s139  (
	.I0(\top/processor/sha_core/n3867_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3867_131 ),
	.I3(\top/processor/sha_core/n3495_171 ),
	.F(\top/processor/sha_core/n3867_115 )
);
defparam \top/processor/sha_core/n3867_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s147  (
	.I0(\top/processor/sha_core/n3607_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [31]),
	.I3(\top/processor/sha_core/w[48] [31]),
	.F(\top/processor/sha_core/n3607_141 )
);
defparam \top/processor/sha_core/n3705_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s147  (
	.I0(\top/processor/sha_core/n3608_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [30]),
	.I3(\top/processor/sha_core/w[48] [30]),
	.F(\top/processor/sha_core/n3608_141 )
);
defparam \top/processor/sha_core/n3706_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s147  (
	.I0(\top/processor/sha_core/n3609_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [29]),
	.I3(\top/processor/sha_core/w[48] [29]),
	.F(\top/processor/sha_core/n3609_141 )
);
defparam \top/processor/sha_core/n3707_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s147  (
	.I0(\top/processor/sha_core/n3610_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [28]),
	.I3(\top/processor/sha_core/w[48] [28]),
	.F(\top/processor/sha_core/n3610_141 )
);
defparam \top/processor/sha_core/n3708_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s147  (
	.I0(\top/processor/sha_core/n3611_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [27]),
	.I3(\top/processor/sha_core/w[48] [27]),
	.F(\top/processor/sha_core/n3611_141 )
);
defparam \top/processor/sha_core/n3709_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s147  (
	.I0(\top/processor/sha_core/n3612_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [26]),
	.I3(\top/processor/sha_core/w[48] [26]),
	.F(\top/processor/sha_core/n3612_141 )
);
defparam \top/processor/sha_core/n3710_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s147  (
	.I0(\top/processor/sha_core/n3613_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [25]),
	.I3(\top/processor/sha_core/w[48] [25]),
	.F(\top/processor/sha_core/n3613_141 )
);
defparam \top/processor/sha_core/n3711_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s147  (
	.I0(\top/processor/sha_core/n3614_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [24]),
	.I3(\top/processor/sha_core/w[48] [24]),
	.F(\top/processor/sha_core/n3614_141 )
);
defparam \top/processor/sha_core/n3712_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s147  (
	.I0(\top/processor/sha_core/n3615_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [23]),
	.I3(\top/processor/sha_core/w[48] [23]),
	.F(\top/processor/sha_core/n3615_141 )
);
defparam \top/processor/sha_core/n3713_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s147  (
	.I0(\top/processor/sha_core/n3616_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [22]),
	.I3(\top/processor/sha_core/w[48] [22]),
	.F(\top/processor/sha_core/n3616_141 )
);
defparam \top/processor/sha_core/n3714_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s147  (
	.I0(\top/processor/sha_core/n3617_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [21]),
	.I3(\top/processor/sha_core/w[48] [21]),
	.F(\top/processor/sha_core/n3617_141 )
);
defparam \top/processor/sha_core/n3715_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s147  (
	.I0(\top/processor/sha_core/n3618_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [20]),
	.I3(\top/processor/sha_core/w[48] [20]),
	.F(\top/processor/sha_core/n3618_141 )
);
defparam \top/processor/sha_core/n3716_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s147  (
	.I0(\top/processor/sha_core/n3619_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [19]),
	.I3(\top/processor/sha_core/w[48] [19]),
	.F(\top/processor/sha_core/n3619_141 )
);
defparam \top/processor/sha_core/n3717_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s147  (
	.I0(\top/processor/sha_core/n3620_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [18]),
	.I3(\top/processor/sha_core/w[48] [18]),
	.F(\top/processor/sha_core/n3620_141 )
);
defparam \top/processor/sha_core/n3718_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s147  (
	.I0(\top/processor/sha_core/n3621_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [17]),
	.I3(\top/processor/sha_core/w[48] [17]),
	.F(\top/processor/sha_core/n3621_141 )
);
defparam \top/processor/sha_core/n3719_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s147  (
	.I0(\top/processor/sha_core/n3622_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [16]),
	.I3(\top/processor/sha_core/w[48] [16]),
	.F(\top/processor/sha_core/n3622_141 )
);
defparam \top/processor/sha_core/n3720_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s147  (
	.I0(\top/processor/sha_core/n3623_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [15]),
	.I3(\top/processor/sha_core/w[48] [15]),
	.F(\top/processor/sha_core/n3623_141 )
);
defparam \top/processor/sha_core/n3721_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s147  (
	.I0(\top/processor/sha_core/n3624_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [14]),
	.I3(\top/processor/sha_core/w[48] [14]),
	.F(\top/processor/sha_core/n3624_141 )
);
defparam \top/processor/sha_core/n3722_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s147  (
	.I0(\top/processor/sha_core/n3625_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [13]),
	.I3(\top/processor/sha_core/w[48] [13]),
	.F(\top/processor/sha_core/n3625_141 )
);
defparam \top/processor/sha_core/n3723_s147 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3496_s180  (
	.I0(\top/processor/sha_core/n3496_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_149 ),
	.I3(\top/processor/sha_core/n3496_150 ),
	.F(\top/processor/sha_core/n3496_133 )
);
defparam \top/processor/sha_core/n3496_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s132  (
	.I0(\top/processor/sha_core/n3868_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_117 ),
	.I3(\top/processor/sha_core/n3496_150 ),
	.F(\top/processor/sha_core/n3868_101 )
);
defparam \top/processor/sha_core/n3868_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3724_s147  (
	.I0(\top/processor/sha_core/n3626_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [12]),
	.I3(\top/processor/sha_core/w[48] [12]),
	.F(\top/processor/sha_core/n3626_141 )
);
defparam \top/processor/sha_core/n3724_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s147  (
	.I0(\top/processor/sha_core/n3627_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [11]),
	.I3(\top/processor/sha_core/w[48] [11]),
	.F(\top/processor/sha_core/n3627_141 )
);
defparam \top/processor/sha_core/n3725_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s147  (
	.I0(\top/processor/sha_core/n3628_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [10]),
	.I3(\top/processor/sha_core/w[48] [10]),
	.F(\top/processor/sha_core/n3628_141 )
);
defparam \top/processor/sha_core/n3726_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s147  (
	.I0(\top/processor/sha_core/n3629_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [9]),
	.I3(\top/processor/sha_core/w[48] [9]),
	.F(\top/processor/sha_core/n3629_141 )
);
defparam \top/processor/sha_core/n3727_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s147  (
	.I0(\top/processor/sha_core/n3630_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [8]),
	.I3(\top/processor/sha_core/w[48] [8]),
	.F(\top/processor/sha_core/n3630_141 )
);
defparam \top/processor/sha_core/n3728_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s147  (
	.I0(\top/processor/sha_core/n3631_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [7]),
	.I3(\top/processor/sha_core/w[48] [7]),
	.F(\top/processor/sha_core/n3631_141 )
);
defparam \top/processor/sha_core/n3729_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s147  (
	.I0(\top/processor/sha_core/n3632_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [6]),
	.I3(\top/processor/sha_core/w[48] [6]),
	.F(\top/processor/sha_core/n3632_141 )
);
defparam \top/processor/sha_core/n3730_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s147  (
	.I0(\top/processor/sha_core/n3633_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [5]),
	.I3(\top/processor/sha_core/w[48] [5]),
	.F(\top/processor/sha_core/n3633_141 )
);
defparam \top/processor/sha_core/n3731_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s147  (
	.I0(\top/processor/sha_core/n3634_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [4]),
	.I3(\top/processor/sha_core/w[48] [4]),
	.F(\top/processor/sha_core/n3634_141 )
);
defparam \top/processor/sha_core/n3732_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s147  (
	.I0(\top/processor/sha_core/n3635_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [3]),
	.I3(\top/processor/sha_core/w[48] [3]),
	.F(\top/processor/sha_core/n3635_141 )
);
defparam \top/processor/sha_core/n3733_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s147  (
	.I0(\top/processor/sha_core/n3636_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [2]),
	.I3(\top/processor/sha_core/w[48] [2]),
	.F(\top/processor/sha_core/n3636_141 )
);
defparam \top/processor/sha_core/n3734_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s147  (
	.I0(\top/processor/sha_core/n3637_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [1]),
	.I3(\top/processor/sha_core/w[48] [1]),
	.F(\top/processor/sha_core/n3637_141 )
);
defparam \top/processor/sha_core/n3735_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s147  (
	.I0(\top/processor/sha_core/n3638_168 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[50] [0]),
	.I3(\top/processor/sha_core/w[48] [0]),
	.F(\top/processor/sha_core/n3638_141 )
);
defparam \top/processor/sha_core/n3736_s147 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3496_s181  (
	.I0(\top/processor/sha_core/n3496_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_152 ),
	.I3(\top/processor/sha_core/n3496_153 ),
	.F(\top/processor/sha_core/n3496_135 )
);
defparam \top/processor/sha_core/n3496_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s133  (
	.I0(\top/processor/sha_core/n3868_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_119 ),
	.I3(\top/processor/sha_core/n3496_153 ),
	.F(\top/processor/sha_core/n3868_103 )
);
defparam \top/processor/sha_core/n3868_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3496_s182  (
	.I0(\top/processor/sha_core/n3496_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_155 ),
	.I3(\top/processor/sha_core/n3496_156 ),
	.F(\top/processor/sha_core/n3496_137 )
);
defparam \top/processor/sha_core/n3496_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s134  (
	.I0(\top/processor/sha_core/n3868_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_121 ),
	.I3(\top/processor/sha_core/n3496_156 ),
	.F(\top/processor/sha_core/n3868_105 )
);
defparam \top/processor/sha_core/n3868_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s148  (
	.I0(\top/processor/sha_core/n3607_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [31]),
	.I3(\top/processor/sha_core/w[52] [31]),
	.F(\top/processor/sha_core/n3607_143 )
);
defparam \top/processor/sha_core/n3705_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s148  (
	.I0(\top/processor/sha_core/n3608_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [30]),
	.I3(\top/processor/sha_core/w[52] [30]),
	.F(\top/processor/sha_core/n3608_143 )
);
defparam \top/processor/sha_core/n3706_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s148  (
	.I0(\top/processor/sha_core/n3609_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [29]),
	.I3(\top/processor/sha_core/w[52] [29]),
	.F(\top/processor/sha_core/n3609_143 )
);
defparam \top/processor/sha_core/n3707_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s148  (
	.I0(\top/processor/sha_core/n3610_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [28]),
	.I3(\top/processor/sha_core/w[52] [28]),
	.F(\top/processor/sha_core/n3610_143 )
);
defparam \top/processor/sha_core/n3708_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s148  (
	.I0(\top/processor/sha_core/n3611_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [27]),
	.I3(\top/processor/sha_core/w[52] [27]),
	.F(\top/processor/sha_core/n3611_143 )
);
defparam \top/processor/sha_core/n3709_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s148  (
	.I0(\top/processor/sha_core/n3612_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [26]),
	.I3(\top/processor/sha_core/w[52] [26]),
	.F(\top/processor/sha_core/n3612_143 )
);
defparam \top/processor/sha_core/n3710_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s148  (
	.I0(\top/processor/sha_core/n3613_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [25]),
	.I3(\top/processor/sha_core/w[52] [25]),
	.F(\top/processor/sha_core/n3613_143 )
);
defparam \top/processor/sha_core/n3711_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s148  (
	.I0(\top/processor/sha_core/n3614_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [24]),
	.I3(\top/processor/sha_core/w[52] [24]),
	.F(\top/processor/sha_core/n3614_143 )
);
defparam \top/processor/sha_core/n3712_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s148  (
	.I0(\top/processor/sha_core/n3615_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [23]),
	.I3(\top/processor/sha_core/w[52] [23]),
	.F(\top/processor/sha_core/n3615_143 )
);
defparam \top/processor/sha_core/n3713_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s148  (
	.I0(\top/processor/sha_core/n3616_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [22]),
	.I3(\top/processor/sha_core/w[52] [22]),
	.F(\top/processor/sha_core/n3616_143 )
);
defparam \top/processor/sha_core/n3714_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s148  (
	.I0(\top/processor/sha_core/n3617_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [21]),
	.I3(\top/processor/sha_core/w[52] [21]),
	.F(\top/processor/sha_core/n3617_143 )
);
defparam \top/processor/sha_core/n3715_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s148  (
	.I0(\top/processor/sha_core/n3618_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [20]),
	.I3(\top/processor/sha_core/w[52] [20]),
	.F(\top/processor/sha_core/n3618_143 )
);
defparam \top/processor/sha_core/n3716_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s148  (
	.I0(\top/processor/sha_core/n3619_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [19]),
	.I3(\top/processor/sha_core/w[52] [19]),
	.F(\top/processor/sha_core/n3619_143 )
);
defparam \top/processor/sha_core/n3717_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s148  (
	.I0(\top/processor/sha_core/n3620_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [18]),
	.I3(\top/processor/sha_core/w[52] [18]),
	.F(\top/processor/sha_core/n3620_143 )
);
defparam \top/processor/sha_core/n3718_s148 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3719_s148  (
	.I0(\top/processor/sha_core/n3621_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [17]),
	.I3(\top/processor/sha_core/w[52] [17]),
	.F(\top/processor/sha_core/n3621_143 )
);
defparam \top/processor/sha_core/n3719_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3496_s183  (
	.I0(\top/processor/sha_core/n3496_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_158 ),
	.I3(\top/processor/sha_core/n3496_159 ),
	.F(\top/processor/sha_core/n3496_139 )
);
defparam \top/processor/sha_core/n3496_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s135  (
	.I0(\top/processor/sha_core/n3868_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_123 ),
	.I3(\top/processor/sha_core/n3496_159 ),
	.F(\top/processor/sha_core/n3868_107 )
);
defparam \top/processor/sha_core/n3868_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3720_s148  (
	.I0(\top/processor/sha_core/n3622_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [16]),
	.I3(\top/processor/sha_core/w[52] [16]),
	.F(\top/processor/sha_core/n3622_143 )
);
defparam \top/processor/sha_core/n3720_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s148  (
	.I0(\top/processor/sha_core/n3623_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [15]),
	.I3(\top/processor/sha_core/w[52] [15]),
	.F(\top/processor/sha_core/n3623_143 )
);
defparam \top/processor/sha_core/n3721_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s148  (
	.I0(\top/processor/sha_core/n3624_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [14]),
	.I3(\top/processor/sha_core/w[52] [14]),
	.F(\top/processor/sha_core/n3624_143 )
);
defparam \top/processor/sha_core/n3722_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s148  (
	.I0(\top/processor/sha_core/n3625_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [13]),
	.I3(\top/processor/sha_core/w[52] [13]),
	.F(\top/processor/sha_core/n3625_143 )
);
defparam \top/processor/sha_core/n3723_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s148  (
	.I0(\top/processor/sha_core/n3626_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [12]),
	.I3(\top/processor/sha_core/w[52] [12]),
	.F(\top/processor/sha_core/n3626_143 )
);
defparam \top/processor/sha_core/n3724_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s148  (
	.I0(\top/processor/sha_core/n3627_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [11]),
	.I3(\top/processor/sha_core/w[52] [11]),
	.F(\top/processor/sha_core/n3627_143 )
);
defparam \top/processor/sha_core/n3725_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s148  (
	.I0(\top/processor/sha_core/n3628_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [10]),
	.I3(\top/processor/sha_core/w[52] [10]),
	.F(\top/processor/sha_core/n3628_143 )
);
defparam \top/processor/sha_core/n3726_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s148  (
	.I0(\top/processor/sha_core/n3629_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [9]),
	.I3(\top/processor/sha_core/w[52] [9]),
	.F(\top/processor/sha_core/n3629_143 )
);
defparam \top/processor/sha_core/n3727_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s148  (
	.I0(\top/processor/sha_core/n3630_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [8]),
	.I3(\top/processor/sha_core/w[52] [8]),
	.F(\top/processor/sha_core/n3630_143 )
);
defparam \top/processor/sha_core/n3728_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s148  (
	.I0(\top/processor/sha_core/n3631_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [7]),
	.I3(\top/processor/sha_core/w[52] [7]),
	.F(\top/processor/sha_core/n3631_143 )
);
defparam \top/processor/sha_core/n3729_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s148  (
	.I0(\top/processor/sha_core/n3632_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [6]),
	.I3(\top/processor/sha_core/w[52] [6]),
	.F(\top/processor/sha_core/n3632_143 )
);
defparam \top/processor/sha_core/n3730_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s148  (
	.I0(\top/processor/sha_core/n3633_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [5]),
	.I3(\top/processor/sha_core/w[52] [5]),
	.F(\top/processor/sha_core/n3633_143 )
);
defparam \top/processor/sha_core/n3731_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s148  (
	.I0(\top/processor/sha_core/n3634_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [4]),
	.I3(\top/processor/sha_core/w[52] [4]),
	.F(\top/processor/sha_core/n3634_143 )
);
defparam \top/processor/sha_core/n3732_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s148  (
	.I0(\top/processor/sha_core/n3635_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [3]),
	.I3(\top/processor/sha_core/w[52] [3]),
	.F(\top/processor/sha_core/n3635_143 )
);
defparam \top/processor/sha_core/n3733_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s148  (
	.I0(\top/processor/sha_core/n3636_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [2]),
	.I3(\top/processor/sha_core/w[52] [2]),
	.F(\top/processor/sha_core/n3636_143 )
);
defparam \top/processor/sha_core/n3734_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s148  (
	.I0(\top/processor/sha_core/n3637_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [1]),
	.I3(\top/processor/sha_core/w[52] [1]),
	.F(\top/processor/sha_core/n3637_143 )
);
defparam \top/processor/sha_core/n3735_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s148  (
	.I0(\top/processor/sha_core/n3638_169 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[54] [0]),
	.I3(\top/processor/sha_core/w[52] [0]),
	.F(\top/processor/sha_core/n3638_143 )
);
defparam \top/processor/sha_core/n3736_s148 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3496_s184  (
	.I0(\top/processor/sha_core/n3496_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_161 ),
	.I3(\top/processor/sha_core/n3496_162 ),
	.F(\top/processor/sha_core/n3496_141 )
);
defparam \top/processor/sha_core/n3496_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s136  (
	.I0(\top/processor/sha_core/n3868_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_125 ),
	.I3(\top/processor/sha_core/n3496_162 ),
	.F(\top/processor/sha_core/n3868_109 )
);
defparam \top/processor/sha_core/n3868_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3496_s185  (
	.I0(\top/processor/sha_core/n3496_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_164 ),
	.I3(\top/processor/sha_core/n3496_165 ),
	.F(\top/processor/sha_core/n3496_143 )
);
defparam \top/processor/sha_core/n3496_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s137  (
	.I0(\top/processor/sha_core/n3868_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_127 ),
	.I3(\top/processor/sha_core/n3496_165 ),
	.F(\top/processor/sha_core/n3868_111 )
);
defparam \top/processor/sha_core/n3868_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s186  (
	.I0(\top/processor/sha_core/n3488_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_152 ),
	.I3(\top/processor/sha_core/n3488_153 ),
	.F(\top/processor/sha_core/n3488_135 )
);
defparam \top/processor/sha_core/n3488_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s138  (
	.I0(\top/processor/sha_core/n3860_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_119 ),
	.I3(\top/processor/sha_core/n3488_153 ),
	.F(\top/processor/sha_core/n3860_103 )
);
defparam \top/processor/sha_core/n3860_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s149  (
	.I0(\top/processor/sha_core/n3607_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [31]),
	.I3(\top/processor/sha_core/w[56] [31]),
	.F(\top/processor/sha_core/n3607_145 )
);
defparam \top/processor/sha_core/n3705_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s149  (
	.I0(\top/processor/sha_core/n3608_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [30]),
	.I3(\top/processor/sha_core/w[56] [30]),
	.F(\top/processor/sha_core/n3608_145 )
);
defparam \top/processor/sha_core/n3706_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s149  (
	.I0(\top/processor/sha_core/n3609_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [29]),
	.I3(\top/processor/sha_core/w[56] [29]),
	.F(\top/processor/sha_core/n3609_145 )
);
defparam \top/processor/sha_core/n3707_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s149  (
	.I0(\top/processor/sha_core/n3610_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [28]),
	.I3(\top/processor/sha_core/w[56] [28]),
	.F(\top/processor/sha_core/n3610_145 )
);
defparam \top/processor/sha_core/n3708_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s149  (
	.I0(\top/processor/sha_core/n3611_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [27]),
	.I3(\top/processor/sha_core/w[56] [27]),
	.F(\top/processor/sha_core/n3611_145 )
);
defparam \top/processor/sha_core/n3709_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s149  (
	.I0(\top/processor/sha_core/n3612_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [26]),
	.I3(\top/processor/sha_core/w[56] [26]),
	.F(\top/processor/sha_core/n3612_145 )
);
defparam \top/processor/sha_core/n3710_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s149  (
	.I0(\top/processor/sha_core/n3613_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [25]),
	.I3(\top/processor/sha_core/w[56] [25]),
	.F(\top/processor/sha_core/n3613_145 )
);
defparam \top/processor/sha_core/n3711_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s149  (
	.I0(\top/processor/sha_core/n3614_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [24]),
	.I3(\top/processor/sha_core/w[56] [24]),
	.F(\top/processor/sha_core/n3614_145 )
);
defparam \top/processor/sha_core/n3712_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s149  (
	.I0(\top/processor/sha_core/n3615_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [23]),
	.I3(\top/processor/sha_core/w[56] [23]),
	.F(\top/processor/sha_core/n3615_145 )
);
defparam \top/processor/sha_core/n3713_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s149  (
	.I0(\top/processor/sha_core/n3616_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [22]),
	.I3(\top/processor/sha_core/w[56] [22]),
	.F(\top/processor/sha_core/n3616_145 )
);
defparam \top/processor/sha_core/n3714_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s149  (
	.I0(\top/processor/sha_core/n3617_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [21]),
	.I3(\top/processor/sha_core/w[56] [21]),
	.F(\top/processor/sha_core/n3617_145 )
);
defparam \top/processor/sha_core/n3715_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3496_s186  (
	.I0(\top/processor/sha_core/n3496_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_167 ),
	.I3(\top/processor/sha_core/n3496_168 ),
	.F(\top/processor/sha_core/n3496_145 )
);
defparam \top/processor/sha_core/n3496_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s138  (
	.I0(\top/processor/sha_core/n3868_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_129 ),
	.I3(\top/processor/sha_core/n3496_168 ),
	.F(\top/processor/sha_core/n3868_113 )
);
defparam \top/processor/sha_core/n3868_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3716_s149  (
	.I0(\top/processor/sha_core/n3618_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [20]),
	.I3(\top/processor/sha_core/w[56] [20]),
	.F(\top/processor/sha_core/n3618_145 )
);
defparam \top/processor/sha_core/n3716_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s149  (
	.I0(\top/processor/sha_core/n3619_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [19]),
	.I3(\top/processor/sha_core/w[56] [19]),
	.F(\top/processor/sha_core/n3619_145 )
);
defparam \top/processor/sha_core/n3717_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s149  (
	.I0(\top/processor/sha_core/n3620_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [18]),
	.I3(\top/processor/sha_core/w[56] [18]),
	.F(\top/processor/sha_core/n3620_145 )
);
defparam \top/processor/sha_core/n3718_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s149  (
	.I0(\top/processor/sha_core/n3621_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [17]),
	.I3(\top/processor/sha_core/w[56] [17]),
	.F(\top/processor/sha_core/n3621_145 )
);
defparam \top/processor/sha_core/n3719_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s149  (
	.I0(\top/processor/sha_core/n3622_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [16]),
	.I3(\top/processor/sha_core/w[56] [16]),
	.F(\top/processor/sha_core/n3622_145 )
);
defparam \top/processor/sha_core/n3720_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s149  (
	.I0(\top/processor/sha_core/n3623_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [15]),
	.I3(\top/processor/sha_core/w[56] [15]),
	.F(\top/processor/sha_core/n3623_145 )
);
defparam \top/processor/sha_core/n3721_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s149  (
	.I0(\top/processor/sha_core/n3624_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [14]),
	.I3(\top/processor/sha_core/w[56] [14]),
	.F(\top/processor/sha_core/n3624_145 )
);
defparam \top/processor/sha_core/n3722_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s149  (
	.I0(\top/processor/sha_core/n3625_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [13]),
	.I3(\top/processor/sha_core/w[56] [13]),
	.F(\top/processor/sha_core/n3625_145 )
);
defparam \top/processor/sha_core/n3723_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s149  (
	.I0(\top/processor/sha_core/n3626_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [12]),
	.I3(\top/processor/sha_core/w[56] [12]),
	.F(\top/processor/sha_core/n3626_145 )
);
defparam \top/processor/sha_core/n3724_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s149  (
	.I0(\top/processor/sha_core/n3627_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [11]),
	.I3(\top/processor/sha_core/w[56] [11]),
	.F(\top/processor/sha_core/n3627_145 )
);
defparam \top/processor/sha_core/n3725_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s149  (
	.I0(\top/processor/sha_core/n3628_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [10]),
	.I3(\top/processor/sha_core/w[56] [10]),
	.F(\top/processor/sha_core/n3628_145 )
);
defparam \top/processor/sha_core/n3726_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s149  (
	.I0(\top/processor/sha_core/n3629_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [9]),
	.I3(\top/processor/sha_core/w[56] [9]),
	.F(\top/processor/sha_core/n3629_145 )
);
defparam \top/processor/sha_core/n3727_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s149  (
	.I0(\top/processor/sha_core/n3630_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [8]),
	.I3(\top/processor/sha_core/w[56] [8]),
	.F(\top/processor/sha_core/n3630_145 )
);
defparam \top/processor/sha_core/n3728_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s149  (
	.I0(\top/processor/sha_core/n3631_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [7]),
	.I3(\top/processor/sha_core/w[56] [7]),
	.F(\top/processor/sha_core/n3631_145 )
);
defparam \top/processor/sha_core/n3729_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s149  (
	.I0(\top/processor/sha_core/n3632_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [6]),
	.I3(\top/processor/sha_core/w[56] [6]),
	.F(\top/processor/sha_core/n3632_145 )
);
defparam \top/processor/sha_core/n3730_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s149  (
	.I0(\top/processor/sha_core/n3633_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [5]),
	.I3(\top/processor/sha_core/w[56] [5]),
	.F(\top/processor/sha_core/n3633_145 )
);
defparam \top/processor/sha_core/n3731_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s149  (
	.I0(\top/processor/sha_core/n3634_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [4]),
	.I3(\top/processor/sha_core/w[56] [4]),
	.F(\top/processor/sha_core/n3634_145 )
);
defparam \top/processor/sha_core/n3732_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s149  (
	.I0(\top/processor/sha_core/n3635_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [3]),
	.I3(\top/processor/sha_core/w[56] [3]),
	.F(\top/processor/sha_core/n3635_145 )
);
defparam \top/processor/sha_core/n3733_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s149  (
	.I0(\top/processor/sha_core/n3636_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [2]),
	.I3(\top/processor/sha_core/w[56] [2]),
	.F(\top/processor/sha_core/n3636_145 )
);
defparam \top/processor/sha_core/n3734_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s149  (
	.I0(\top/processor/sha_core/n3637_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [1]),
	.I3(\top/processor/sha_core/w[56] [1]),
	.F(\top/processor/sha_core/n3637_145 )
);
defparam \top/processor/sha_core/n3735_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3496_s187  (
	.I0(\top/processor/sha_core/n3496_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_170 ),
	.I3(\top/processor/sha_core/n3496_171 ),
	.F(\top/processor/sha_core/n3496_147 )
);
defparam \top/processor/sha_core/n3496_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3868_s139  (
	.I0(\top/processor/sha_core/n3868_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3868_131 ),
	.I3(\top/processor/sha_core/n3496_171 ),
	.F(\top/processor/sha_core/n3868_115 )
);
defparam \top/processor/sha_core/n3868_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3736_s149  (
	.I0(\top/processor/sha_core/n3638_170 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[58] [0]),
	.I3(\top/processor/sha_core/w[56] [0]),
	.F(\top/processor/sha_core/n3638_145 )
);
defparam \top/processor/sha_core/n3736_s149 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3497_s180  (
	.I0(\top/processor/sha_core/n3497_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_149 ),
	.I3(\top/processor/sha_core/n3497_150 ),
	.F(\top/processor/sha_core/n3497_133 )
);
defparam \top/processor/sha_core/n3497_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s132  (
	.I0(\top/processor/sha_core/n3869_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_117 ),
	.I3(\top/processor/sha_core/n3497_150 ),
	.F(\top/processor/sha_core/n3869_101 )
);
defparam \top/processor/sha_core/n3869_s132 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3705_s150  (
	.I0(\top/processor/sha_core/n3607_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [31]),
	.I3(\top/processor/sha_core/w[60] [31]),
	.F(\top/processor/sha_core/n3607_147 )
);
defparam \top/processor/sha_core/n3705_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s150  (
	.I0(\top/processor/sha_core/n3608_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [30]),
	.I3(\top/processor/sha_core/w[60] [30]),
	.F(\top/processor/sha_core/n3608_147 )
);
defparam \top/processor/sha_core/n3706_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s150  (
	.I0(\top/processor/sha_core/n3609_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [29]),
	.I3(\top/processor/sha_core/w[60] [29]),
	.F(\top/processor/sha_core/n3609_147 )
);
defparam \top/processor/sha_core/n3707_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s150  (
	.I0(\top/processor/sha_core/n3610_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [28]),
	.I3(\top/processor/sha_core/w[60] [28]),
	.F(\top/processor/sha_core/n3610_147 )
);
defparam \top/processor/sha_core/n3708_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s150  (
	.I0(\top/processor/sha_core/n3611_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [27]),
	.I3(\top/processor/sha_core/w[60] [27]),
	.F(\top/processor/sha_core/n3611_147 )
);
defparam \top/processor/sha_core/n3709_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s150  (
	.I0(\top/processor/sha_core/n3612_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [26]),
	.I3(\top/processor/sha_core/w[60] [26]),
	.F(\top/processor/sha_core/n3612_147 )
);
defparam \top/processor/sha_core/n3710_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s150  (
	.I0(\top/processor/sha_core/n3613_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [25]),
	.I3(\top/processor/sha_core/w[60] [25]),
	.F(\top/processor/sha_core/n3613_147 )
);
defparam \top/processor/sha_core/n3711_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3497_s181  (
	.I0(\top/processor/sha_core/n3497_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_152 ),
	.I3(\top/processor/sha_core/n3497_153 ),
	.F(\top/processor/sha_core/n3497_135 )
);
defparam \top/processor/sha_core/n3497_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s133  (
	.I0(\top/processor/sha_core/n3869_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_119 ),
	.I3(\top/processor/sha_core/n3497_153 ),
	.F(\top/processor/sha_core/n3869_103 )
);
defparam \top/processor/sha_core/n3869_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3712_s150  (
	.I0(\top/processor/sha_core/n3614_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [24]),
	.I3(\top/processor/sha_core/w[60] [24]),
	.F(\top/processor/sha_core/n3614_147 )
);
defparam \top/processor/sha_core/n3712_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s150  (
	.I0(\top/processor/sha_core/n3615_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [23]),
	.I3(\top/processor/sha_core/w[60] [23]),
	.F(\top/processor/sha_core/n3615_147 )
);
defparam \top/processor/sha_core/n3713_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s150  (
	.I0(\top/processor/sha_core/n3616_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [22]),
	.I3(\top/processor/sha_core/w[60] [22]),
	.F(\top/processor/sha_core/n3616_147 )
);
defparam \top/processor/sha_core/n3714_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s150  (
	.I0(\top/processor/sha_core/n3617_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [21]),
	.I3(\top/processor/sha_core/w[60] [21]),
	.F(\top/processor/sha_core/n3617_147 )
);
defparam \top/processor/sha_core/n3715_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s150  (
	.I0(\top/processor/sha_core/n3618_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [20]),
	.I3(\top/processor/sha_core/w[60] [20]),
	.F(\top/processor/sha_core/n3618_147 )
);
defparam \top/processor/sha_core/n3716_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s150  (
	.I0(\top/processor/sha_core/n3619_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [19]),
	.I3(\top/processor/sha_core/w[60] [19]),
	.F(\top/processor/sha_core/n3619_147 )
);
defparam \top/processor/sha_core/n3717_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s150  (
	.I0(\top/processor/sha_core/n3620_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [18]),
	.I3(\top/processor/sha_core/w[60] [18]),
	.F(\top/processor/sha_core/n3620_147 )
);
defparam \top/processor/sha_core/n3718_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s150  (
	.I0(\top/processor/sha_core/n3621_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [17]),
	.I3(\top/processor/sha_core/w[60] [17]),
	.F(\top/processor/sha_core/n3621_147 )
);
defparam \top/processor/sha_core/n3719_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s150  (
	.I0(\top/processor/sha_core/n3622_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [16]),
	.I3(\top/processor/sha_core/w[60] [16]),
	.F(\top/processor/sha_core/n3622_147 )
);
defparam \top/processor/sha_core/n3720_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s150  (
	.I0(\top/processor/sha_core/n3623_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [15]),
	.I3(\top/processor/sha_core/w[60] [15]),
	.F(\top/processor/sha_core/n3623_147 )
);
defparam \top/processor/sha_core/n3721_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s150  (
	.I0(\top/processor/sha_core/n3624_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [14]),
	.I3(\top/processor/sha_core/w[60] [14]),
	.F(\top/processor/sha_core/n3624_147 )
);
defparam \top/processor/sha_core/n3722_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s150  (
	.I0(\top/processor/sha_core/n3625_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [13]),
	.I3(\top/processor/sha_core/w[60] [13]),
	.F(\top/processor/sha_core/n3625_147 )
);
defparam \top/processor/sha_core/n3723_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s150  (
	.I0(\top/processor/sha_core/n3626_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [12]),
	.I3(\top/processor/sha_core/w[60] [12]),
	.F(\top/processor/sha_core/n3626_147 )
);
defparam \top/processor/sha_core/n3724_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s150  (
	.I0(\top/processor/sha_core/n3627_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [11]),
	.I3(\top/processor/sha_core/w[60] [11]),
	.F(\top/processor/sha_core/n3627_147 )
);
defparam \top/processor/sha_core/n3725_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s150  (
	.I0(\top/processor/sha_core/n3628_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [10]),
	.I3(\top/processor/sha_core/w[60] [10]),
	.F(\top/processor/sha_core/n3628_147 )
);
defparam \top/processor/sha_core/n3726_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s150  (
	.I0(\top/processor/sha_core/n3629_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [9]),
	.I3(\top/processor/sha_core/w[60] [9]),
	.F(\top/processor/sha_core/n3629_147 )
);
defparam \top/processor/sha_core/n3727_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s150  (
	.I0(\top/processor/sha_core/n3630_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [8]),
	.I3(\top/processor/sha_core/w[60] [8]),
	.F(\top/processor/sha_core/n3630_147 )
);
defparam \top/processor/sha_core/n3728_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s150  (
	.I0(\top/processor/sha_core/n3631_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [7]),
	.I3(\top/processor/sha_core/w[60] [7]),
	.F(\top/processor/sha_core/n3631_147 )
);
defparam \top/processor/sha_core/n3729_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s150  (
	.I0(\top/processor/sha_core/n3632_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [6]),
	.I3(\top/processor/sha_core/w[60] [6]),
	.F(\top/processor/sha_core/n3632_147 )
);
defparam \top/processor/sha_core/n3730_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s150  (
	.I0(\top/processor/sha_core/n3633_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [5]),
	.I3(\top/processor/sha_core/w[60] [5]),
	.F(\top/processor/sha_core/n3633_147 )
);
defparam \top/processor/sha_core/n3731_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3497_s182  (
	.I0(\top/processor/sha_core/n3497_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_155 ),
	.I3(\top/processor/sha_core/n3497_156 ),
	.F(\top/processor/sha_core/n3497_137 )
);
defparam \top/processor/sha_core/n3497_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s134  (
	.I0(\top/processor/sha_core/n3869_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_121 ),
	.I3(\top/processor/sha_core/n3497_156 ),
	.F(\top/processor/sha_core/n3869_105 )
);
defparam \top/processor/sha_core/n3869_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3732_s150  (
	.I0(\top/processor/sha_core/n3634_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [4]),
	.I3(\top/processor/sha_core/w[60] [4]),
	.F(\top/processor/sha_core/n3634_147 )
);
defparam \top/processor/sha_core/n3732_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s150  (
	.I0(\top/processor/sha_core/n3635_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [3]),
	.I3(\top/processor/sha_core/w[60] [3]),
	.F(\top/processor/sha_core/n3635_147 )
);
defparam \top/processor/sha_core/n3733_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s150  (
	.I0(\top/processor/sha_core/n3636_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [2]),
	.I3(\top/processor/sha_core/w[60] [2]),
	.F(\top/processor/sha_core/n3636_147 )
);
defparam \top/processor/sha_core/n3734_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s150  (
	.I0(\top/processor/sha_core/n3637_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [1]),
	.I3(\top/processor/sha_core/w[60] [1]),
	.F(\top/processor/sha_core/n3637_147 )
);
defparam \top/processor/sha_core/n3735_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s150  (
	.I0(\top/processor/sha_core/n3638_171 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[62] [0]),
	.I3(\top/processor/sha_core/w[60] [0]),
	.F(\top/processor/sha_core/n3638_147 )
);
defparam \top/processor/sha_core/n3736_s150 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3497_s183  (
	.I0(\top/processor/sha_core/n3497_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_158 ),
	.I3(\top/processor/sha_core/n3497_159 ),
	.F(\top/processor/sha_core/n3497_139 )
);
defparam \top/processor/sha_core/n3497_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s135  (
	.I0(\top/processor/sha_core/n3869_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_123 ),
	.I3(\top/processor/sha_core/n3497_159 ),
	.F(\top/processor/sha_core/n3869_107 )
);
defparam \top/processor/sha_core/n3869_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3497_s184  (
	.I0(\top/processor/sha_core/n3497_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_161 ),
	.I3(\top/processor/sha_core/n3497_162 ),
	.F(\top/processor/sha_core/n3497_141 )
);
defparam \top/processor/sha_core/n3497_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s136  (
	.I0(\top/processor/sha_core/n3869_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_125 ),
	.I3(\top/processor/sha_core/n3497_162 ),
	.F(\top/processor/sha_core/n3869_109 )
);
defparam \top/processor/sha_core/n3869_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3497_s185  (
	.I0(\top/processor/sha_core/n3497_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_164 ),
	.I3(\top/processor/sha_core/n3497_165 ),
	.F(\top/processor/sha_core/n3497_143 )
);
defparam \top/processor/sha_core/n3497_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s137  (
	.I0(\top/processor/sha_core/n3869_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_127 ),
	.I3(\top/processor/sha_core/n3497_165 ),
	.F(\top/processor/sha_core/n3869_111 )
);
defparam \top/processor/sha_core/n3869_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3497_s186  (
	.I0(\top/processor/sha_core/n3497_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_167 ),
	.I3(\top/processor/sha_core/n3497_168 ),
	.F(\top/processor/sha_core/n3497_145 )
);
defparam \top/processor/sha_core/n3497_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s138  (
	.I0(\top/processor/sha_core/n3869_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_129 ),
	.I3(\top/processor/sha_core/n3497_168 ),
	.F(\top/processor/sha_core/n3869_113 )
);
defparam \top/processor/sha_core/n3869_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3497_s187  (
	.I0(\top/processor/sha_core/n3497_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_170 ),
	.I3(\top/processor/sha_core/n3497_171 ),
	.F(\top/processor/sha_core/n3497_147 )
);
defparam \top/processor/sha_core/n3497_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3869_s139  (
	.I0(\top/processor/sha_core/n3869_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3869_131 ),
	.I3(\top/processor/sha_core/n3497_171 ),
	.F(\top/processor/sha_core/n3869_115 )
);
defparam \top/processor/sha_core/n3869_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s187  (
	.I0(\top/processor/sha_core/n3488_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_155 ),
	.I3(\top/processor/sha_core/n3488_156 ),
	.F(\top/processor/sha_core/n3488_137 )
);
defparam \top/processor/sha_core/n3488_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s139  (
	.I0(\top/processor/sha_core/n3860_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_121 ),
	.I3(\top/processor/sha_core/n3488_156 ),
	.F(\top/processor/sha_core/n3860_105 )
);
defparam \top/processor/sha_core/n3860_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s180  (
	.I0(\top/processor/sha_core/n3498_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_149 ),
	.I3(\top/processor/sha_core/n3498_150 ),
	.F(\top/processor/sha_core/n3498_133 )
);
defparam \top/processor/sha_core/n3498_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s132  (
	.I0(\top/processor/sha_core/n3870_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_117 ),
	.I3(\top/processor/sha_core/n3498_150 ),
	.F(\top/processor/sha_core/n3870_101 )
);
defparam \top/processor/sha_core/n3870_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s181  (
	.I0(\top/processor/sha_core/n3498_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_152 ),
	.I3(\top/processor/sha_core/n3498_153 ),
	.F(\top/processor/sha_core/n3498_135 )
);
defparam \top/processor/sha_core/n3498_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s133  (
	.I0(\top/processor/sha_core/n3870_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_119 ),
	.I3(\top/processor/sha_core/n3498_153 ),
	.F(\top/processor/sha_core/n3870_103 )
);
defparam \top/processor/sha_core/n3870_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s182  (
	.I0(\top/processor/sha_core/n3498_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_155 ),
	.I3(\top/processor/sha_core/n3498_156 ),
	.F(\top/processor/sha_core/n3498_137 )
);
defparam \top/processor/sha_core/n3498_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s134  (
	.I0(\top/processor/sha_core/n3870_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_121 ),
	.I3(\top/processor/sha_core/n3498_156 ),
	.F(\top/processor/sha_core/n3870_105 )
);
defparam \top/processor/sha_core/n3870_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s183  (
	.I0(\top/processor/sha_core/n3498_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_158 ),
	.I3(\top/processor/sha_core/n3498_159 ),
	.F(\top/processor/sha_core/n3498_139 )
);
defparam \top/processor/sha_core/n3498_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s135  (
	.I0(\top/processor/sha_core/n3870_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_123 ),
	.I3(\top/processor/sha_core/n3498_159 ),
	.F(\top/processor/sha_core/n3870_107 )
);
defparam \top/processor/sha_core/n3870_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s184  (
	.I0(\top/processor/sha_core/n3498_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_161 ),
	.I3(\top/processor/sha_core/n3498_162 ),
	.F(\top/processor/sha_core/n3498_141 )
);
defparam \top/processor/sha_core/n3498_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s136  (
	.I0(\top/processor/sha_core/n3870_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_125 ),
	.I3(\top/processor/sha_core/n3498_162 ),
	.F(\top/processor/sha_core/n3870_109 )
);
defparam \top/processor/sha_core/n3870_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s185  (
	.I0(\top/processor/sha_core/n3498_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_164 ),
	.I3(\top/processor/sha_core/n3498_165 ),
	.F(\top/processor/sha_core/n3498_143 )
);
defparam \top/processor/sha_core/n3498_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s137  (
	.I0(\top/processor/sha_core/n3870_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_127 ),
	.I3(\top/processor/sha_core/n3498_165 ),
	.F(\top/processor/sha_core/n3870_111 )
);
defparam \top/processor/sha_core/n3870_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s186  (
	.I0(\top/processor/sha_core/n3498_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_167 ),
	.I3(\top/processor/sha_core/n3498_168 ),
	.F(\top/processor/sha_core/n3498_145 )
);
defparam \top/processor/sha_core/n3498_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s138  (
	.I0(\top/processor/sha_core/n3870_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_129 ),
	.I3(\top/processor/sha_core/n3498_168 ),
	.F(\top/processor/sha_core/n3870_113 )
);
defparam \top/processor/sha_core/n3870_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3498_s187  (
	.I0(\top/processor/sha_core/n3498_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_170 ),
	.I3(\top/processor/sha_core/n3498_171 ),
	.F(\top/processor/sha_core/n3498_147 )
);
defparam \top/processor/sha_core/n3498_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3870_s139  (
	.I0(\top/processor/sha_core/n3870_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3870_131 ),
	.I3(\top/processor/sha_core/n3498_171 ),
	.F(\top/processor/sha_core/n3870_115 )
);
defparam \top/processor/sha_core/n3870_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s180  (
	.I0(\top/processor/sha_core/n3499_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_149 ),
	.I3(\top/processor/sha_core/n3499_150 ),
	.F(\top/processor/sha_core/n3499_133 )
);
defparam \top/processor/sha_core/n3499_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s132  (
	.I0(\top/processor/sha_core/n3871_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_117 ),
	.I3(\top/processor/sha_core/n3499_150 ),
	.F(\top/processor/sha_core/n3871_101 )
);
defparam \top/processor/sha_core/n3871_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s181  (
	.I0(\top/processor/sha_core/n3499_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_152 ),
	.I3(\top/processor/sha_core/n3499_153 ),
	.F(\top/processor/sha_core/n3499_135 )
);
defparam \top/processor/sha_core/n3499_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s133  (
	.I0(\top/processor/sha_core/n3871_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_119 ),
	.I3(\top/processor/sha_core/n3499_153 ),
	.F(\top/processor/sha_core/n3871_103 )
);
defparam \top/processor/sha_core/n3871_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s180  (
	.I0(\top/processor/sha_core/n3489_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_149 ),
	.I3(\top/processor/sha_core/n3489_150 ),
	.F(\top/processor/sha_core/n3489_133 )
);
defparam \top/processor/sha_core/n3489_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s132  (
	.I0(\top/processor/sha_core/n3861_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_117 ),
	.I3(\top/processor/sha_core/n3489_150 ),
	.F(\top/processor/sha_core/n3861_101 )
);
defparam \top/processor/sha_core/n3861_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s182  (
	.I0(\top/processor/sha_core/n3499_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_155 ),
	.I3(\top/processor/sha_core/n3499_156 ),
	.F(\top/processor/sha_core/n3499_137 )
);
defparam \top/processor/sha_core/n3499_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s134  (
	.I0(\top/processor/sha_core/n3871_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_121 ),
	.I3(\top/processor/sha_core/n3499_156 ),
	.F(\top/processor/sha_core/n3871_105 )
);
defparam \top/processor/sha_core/n3871_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s183  (
	.I0(\top/processor/sha_core/n3499_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_158 ),
	.I3(\top/processor/sha_core/n3499_159 ),
	.F(\top/processor/sha_core/n3499_139 )
);
defparam \top/processor/sha_core/n3499_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s135  (
	.I0(\top/processor/sha_core/n3871_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_123 ),
	.I3(\top/processor/sha_core/n3499_159 ),
	.F(\top/processor/sha_core/n3871_107 )
);
defparam \top/processor/sha_core/n3871_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s184  (
	.I0(\top/processor/sha_core/n3499_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_161 ),
	.I3(\top/processor/sha_core/n3499_162 ),
	.F(\top/processor/sha_core/n3499_141 )
);
defparam \top/processor/sha_core/n3499_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s136  (
	.I0(\top/processor/sha_core/n3871_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_125 ),
	.I3(\top/processor/sha_core/n3499_162 ),
	.F(\top/processor/sha_core/n3871_109 )
);
defparam \top/processor/sha_core/n3871_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s185  (
	.I0(\top/processor/sha_core/n3499_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_164 ),
	.I3(\top/processor/sha_core/n3499_165 ),
	.F(\top/processor/sha_core/n3499_143 )
);
defparam \top/processor/sha_core/n3499_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s137  (
	.I0(\top/processor/sha_core/n3871_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_127 ),
	.I3(\top/processor/sha_core/n3499_165 ),
	.F(\top/processor/sha_core/n3871_111 )
);
defparam \top/processor/sha_core/n3871_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s186  (
	.I0(\top/processor/sha_core/n3499_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_167 ),
	.I3(\top/processor/sha_core/n3499_168 ),
	.F(\top/processor/sha_core/n3499_145 )
);
defparam \top/processor/sha_core/n3499_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s138  (
	.I0(\top/processor/sha_core/n3871_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_129 ),
	.I3(\top/processor/sha_core/n3499_168 ),
	.F(\top/processor/sha_core/n3871_113 )
);
defparam \top/processor/sha_core/n3871_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3499_s187  (
	.I0(\top/processor/sha_core/n3499_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_170 ),
	.I3(\top/processor/sha_core/n3499_171 ),
	.F(\top/processor/sha_core/n3499_147 )
);
defparam \top/processor/sha_core/n3499_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3871_s139  (
	.I0(\top/processor/sha_core/n3871_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3871_131 ),
	.I3(\top/processor/sha_core/n3499_171 ),
	.F(\top/processor/sha_core/n3871_115 )
);
defparam \top/processor/sha_core/n3871_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s180  (
	.I0(\top/processor/sha_core/n3500_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_149 ),
	.I3(\top/processor/sha_core/n3500_150 ),
	.F(\top/processor/sha_core/n3500_133 )
);
defparam \top/processor/sha_core/n3500_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s132  (
	.I0(\top/processor/sha_core/n3872_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_117 ),
	.I3(\top/processor/sha_core/n3500_150 ),
	.F(\top/processor/sha_core/n3872_101 )
);
defparam \top/processor/sha_core/n3872_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s181  (
	.I0(\top/processor/sha_core/n3500_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_152 ),
	.I3(\top/processor/sha_core/n3500_153 ),
	.F(\top/processor/sha_core/n3500_135 )
);
defparam \top/processor/sha_core/n3500_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s133  (
	.I0(\top/processor/sha_core/n3872_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_119 ),
	.I3(\top/processor/sha_core/n3500_153 ),
	.F(\top/processor/sha_core/n3872_103 )
);
defparam \top/processor/sha_core/n3872_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s182  (
	.I0(\top/processor/sha_core/n3500_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_155 ),
	.I3(\top/processor/sha_core/n3500_156 ),
	.F(\top/processor/sha_core/n3500_137 )
);
defparam \top/processor/sha_core/n3500_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s134  (
	.I0(\top/processor/sha_core/n3872_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_121 ),
	.I3(\top/processor/sha_core/n3500_156 ),
	.F(\top/processor/sha_core/n3872_105 )
);
defparam \top/processor/sha_core/n3872_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s183  (
	.I0(\top/processor/sha_core/n3500_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_158 ),
	.I3(\top/processor/sha_core/n3500_159 ),
	.F(\top/processor/sha_core/n3500_139 )
);
defparam \top/processor/sha_core/n3500_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s135  (
	.I0(\top/processor/sha_core/n3872_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_123 ),
	.I3(\top/processor/sha_core/n3500_159 ),
	.F(\top/processor/sha_core/n3872_107 )
);
defparam \top/processor/sha_core/n3872_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s181  (
	.I0(\top/processor/sha_core/n3489_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_152 ),
	.I3(\top/processor/sha_core/n3489_153 ),
	.F(\top/processor/sha_core/n3489_135 )
);
defparam \top/processor/sha_core/n3489_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s133  (
	.I0(\top/processor/sha_core/n3861_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_119 ),
	.I3(\top/processor/sha_core/n3489_153 ),
	.F(\top/processor/sha_core/n3861_103 )
);
defparam \top/processor/sha_core/n3861_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s180  (
	.I0(\top/processor/sha_core/n3488_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_158 ),
	.I3(\top/processor/sha_core/n3488_159 ),
	.F(\top/processor/sha_core/n3488_139 )
);
defparam \top/processor/sha_core/n3488_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s132  (
	.I0(\top/processor/sha_core/n3860_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_123 ),
	.I3(\top/processor/sha_core/n3488_159 ),
	.F(\top/processor/sha_core/n3860_107 )
);
defparam \top/processor/sha_core/n3860_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s184  (
	.I0(\top/processor/sha_core/n3500_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_161 ),
	.I3(\top/processor/sha_core/n3500_162 ),
	.F(\top/processor/sha_core/n3500_141 )
);
defparam \top/processor/sha_core/n3500_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s136  (
	.I0(\top/processor/sha_core/n3872_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_125 ),
	.I3(\top/processor/sha_core/n3500_162 ),
	.F(\top/processor/sha_core/n3872_109 )
);
defparam \top/processor/sha_core/n3872_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s185  (
	.I0(\top/processor/sha_core/n3500_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_164 ),
	.I3(\top/processor/sha_core/n3500_165 ),
	.F(\top/processor/sha_core/n3500_143 )
);
defparam \top/processor/sha_core/n3500_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s137  (
	.I0(\top/processor/sha_core/n3872_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_127 ),
	.I3(\top/processor/sha_core/n3500_165 ),
	.F(\top/processor/sha_core/n3872_111 )
);
defparam \top/processor/sha_core/n3872_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s186  (
	.I0(\top/processor/sha_core/n3500_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_167 ),
	.I3(\top/processor/sha_core/n3500_168 ),
	.F(\top/processor/sha_core/n3500_145 )
);
defparam \top/processor/sha_core/n3500_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s138  (
	.I0(\top/processor/sha_core/n3872_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_129 ),
	.I3(\top/processor/sha_core/n3500_168 ),
	.F(\top/processor/sha_core/n3872_113 )
);
defparam \top/processor/sha_core/n3872_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3500_s187  (
	.I0(\top/processor/sha_core/n3500_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_170 ),
	.I3(\top/processor/sha_core/n3500_171 ),
	.F(\top/processor/sha_core/n3500_147 )
);
defparam \top/processor/sha_core/n3500_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3872_s139  (
	.I0(\top/processor/sha_core/n3872_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3872_131 ),
	.I3(\top/processor/sha_core/n3500_171 ),
	.F(\top/processor/sha_core/n3872_115 )
);
defparam \top/processor/sha_core/n3872_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s180  (
	.I0(\top/processor/sha_core/n3501_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_149 ),
	.I3(\top/processor/sha_core/n3501_150 ),
	.F(\top/processor/sha_core/n3501_133 )
);
defparam \top/processor/sha_core/n3501_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s132  (
	.I0(\top/processor/sha_core/n3873_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_117 ),
	.I3(\top/processor/sha_core/n3501_150 ),
	.F(\top/processor/sha_core/n3873_101 )
);
defparam \top/processor/sha_core/n3873_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s181  (
	.I0(\top/processor/sha_core/n3501_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_152 ),
	.I3(\top/processor/sha_core/n3501_153 ),
	.F(\top/processor/sha_core/n3501_135 )
);
defparam \top/processor/sha_core/n3501_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s133  (
	.I0(\top/processor/sha_core/n3873_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_119 ),
	.I3(\top/processor/sha_core/n3501_153 ),
	.F(\top/processor/sha_core/n3873_103 )
);
defparam \top/processor/sha_core/n3873_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s182  (
	.I0(\top/processor/sha_core/n3501_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_155 ),
	.I3(\top/processor/sha_core/n3501_156 ),
	.F(\top/processor/sha_core/n3501_137 )
);
defparam \top/processor/sha_core/n3501_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s134  (
	.I0(\top/processor/sha_core/n3873_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_121 ),
	.I3(\top/processor/sha_core/n3501_156 ),
	.F(\top/processor/sha_core/n3873_105 )
);
defparam \top/processor/sha_core/n3873_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s183  (
	.I0(\top/processor/sha_core/n3501_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_158 ),
	.I3(\top/processor/sha_core/n3501_159 ),
	.F(\top/processor/sha_core/n3501_139 )
);
defparam \top/processor/sha_core/n3501_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s135  (
	.I0(\top/processor/sha_core/n3873_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_123 ),
	.I3(\top/processor/sha_core/n3501_159 ),
	.F(\top/processor/sha_core/n3873_107 )
);
defparam \top/processor/sha_core/n3873_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s184  (
	.I0(\top/processor/sha_core/n3501_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_161 ),
	.I3(\top/processor/sha_core/n3501_162 ),
	.F(\top/processor/sha_core/n3501_141 )
);
defparam \top/processor/sha_core/n3501_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s136  (
	.I0(\top/processor/sha_core/n3873_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_125 ),
	.I3(\top/processor/sha_core/n3501_162 ),
	.F(\top/processor/sha_core/n3873_109 )
);
defparam \top/processor/sha_core/n3873_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s185  (
	.I0(\top/processor/sha_core/n3501_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_164 ),
	.I3(\top/processor/sha_core/n3501_165 ),
	.F(\top/processor/sha_core/n3501_143 )
);
defparam \top/processor/sha_core/n3501_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s137  (
	.I0(\top/processor/sha_core/n3873_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_127 ),
	.I3(\top/processor/sha_core/n3501_165 ),
	.F(\top/processor/sha_core/n3873_111 )
);
defparam \top/processor/sha_core/n3873_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s182  (
	.I0(\top/processor/sha_core/n3489_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_155 ),
	.I3(\top/processor/sha_core/n3489_156 ),
	.F(\top/processor/sha_core/n3489_137 )
);
defparam \top/processor/sha_core/n3489_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s134  (
	.I0(\top/processor/sha_core/n3861_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_121 ),
	.I3(\top/processor/sha_core/n3489_156 ),
	.F(\top/processor/sha_core/n3861_105 )
);
defparam \top/processor/sha_core/n3861_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s186  (
	.I0(\top/processor/sha_core/n3501_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_167 ),
	.I3(\top/processor/sha_core/n3501_168 ),
	.F(\top/processor/sha_core/n3501_145 )
);
defparam \top/processor/sha_core/n3501_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s138  (
	.I0(\top/processor/sha_core/n3873_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_129 ),
	.I3(\top/processor/sha_core/n3501_168 ),
	.F(\top/processor/sha_core/n3873_113 )
);
defparam \top/processor/sha_core/n3873_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3501_s187  (
	.I0(\top/processor/sha_core/n3501_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_170 ),
	.I3(\top/processor/sha_core/n3501_171 ),
	.F(\top/processor/sha_core/n3501_147 )
);
defparam \top/processor/sha_core/n3501_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3873_s139  (
	.I0(\top/processor/sha_core/n3873_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3873_131 ),
	.I3(\top/processor/sha_core/n3501_171 ),
	.F(\top/processor/sha_core/n3873_115 )
);
defparam \top/processor/sha_core/n3873_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s180  (
	.I0(\top/processor/sha_core/n3502_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_149 ),
	.I3(\top/processor/sha_core/n3502_150 ),
	.F(\top/processor/sha_core/n3502_133 )
);
defparam \top/processor/sha_core/n3502_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s132  (
	.I0(\top/processor/sha_core/n3874_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_117 ),
	.I3(\top/processor/sha_core/n3502_150 ),
	.F(\top/processor/sha_core/n3874_101 )
);
defparam \top/processor/sha_core/n3874_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s181  (
	.I0(\top/processor/sha_core/n3502_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_152 ),
	.I3(\top/processor/sha_core/n3502_153 ),
	.F(\top/processor/sha_core/n3502_135 )
);
defparam \top/processor/sha_core/n3502_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s133  (
	.I0(\top/processor/sha_core/n3874_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_119 ),
	.I3(\top/processor/sha_core/n3502_153 ),
	.F(\top/processor/sha_core/n3874_103 )
);
defparam \top/processor/sha_core/n3874_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s182  (
	.I0(\top/processor/sha_core/n3502_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_155 ),
	.I3(\top/processor/sha_core/n3502_156 ),
	.F(\top/processor/sha_core/n3502_137 )
);
defparam \top/processor/sha_core/n3502_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s134  (
	.I0(\top/processor/sha_core/n3874_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_121 ),
	.I3(\top/processor/sha_core/n3502_156 ),
	.F(\top/processor/sha_core/n3874_105 )
);
defparam \top/processor/sha_core/n3874_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s183  (
	.I0(\top/processor/sha_core/n3502_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_158 ),
	.I3(\top/processor/sha_core/n3502_159 ),
	.F(\top/processor/sha_core/n3502_139 )
);
defparam \top/processor/sha_core/n3502_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s135  (
	.I0(\top/processor/sha_core/n3874_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_123 ),
	.I3(\top/processor/sha_core/n3502_159 ),
	.F(\top/processor/sha_core/n3874_107 )
);
defparam \top/processor/sha_core/n3874_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s184  (
	.I0(\top/processor/sha_core/n3502_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_161 ),
	.I3(\top/processor/sha_core/n3502_162 ),
	.F(\top/processor/sha_core/n3502_141 )
);
defparam \top/processor/sha_core/n3502_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s136  (
	.I0(\top/processor/sha_core/n3874_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_125 ),
	.I3(\top/processor/sha_core/n3502_162 ),
	.F(\top/processor/sha_core/n3874_109 )
);
defparam \top/processor/sha_core/n3874_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s185  (
	.I0(\top/processor/sha_core/n3502_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_164 ),
	.I3(\top/processor/sha_core/n3502_165 ),
	.F(\top/processor/sha_core/n3502_143 )
);
defparam \top/processor/sha_core/n3502_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s137  (
	.I0(\top/processor/sha_core/n3874_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_127 ),
	.I3(\top/processor/sha_core/n3502_165 ),
	.F(\top/processor/sha_core/n3874_111 )
);
defparam \top/processor/sha_core/n3874_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s186  (
	.I0(\top/processor/sha_core/n3502_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_167 ),
	.I3(\top/processor/sha_core/n3502_168 ),
	.F(\top/processor/sha_core/n3502_145 )
);
defparam \top/processor/sha_core/n3502_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s138  (
	.I0(\top/processor/sha_core/n3874_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_129 ),
	.I3(\top/processor/sha_core/n3502_168 ),
	.F(\top/processor/sha_core/n3874_113 )
);
defparam \top/processor/sha_core/n3874_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3502_s187  (
	.I0(\top/processor/sha_core/n3502_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_170 ),
	.I3(\top/processor/sha_core/n3502_171 ),
	.F(\top/processor/sha_core/n3502_147 )
);
defparam \top/processor/sha_core/n3502_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3874_s139  (
	.I0(\top/processor/sha_core/n3874_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3874_131 ),
	.I3(\top/processor/sha_core/n3502_171 ),
	.F(\top/processor/sha_core/n3874_115 )
);
defparam \top/processor/sha_core/n3874_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s183  (
	.I0(\top/processor/sha_core/n3489_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_158 ),
	.I3(\top/processor/sha_core/n3489_159 ),
	.F(\top/processor/sha_core/n3489_139 )
);
defparam \top/processor/sha_core/n3489_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s135  (
	.I0(\top/processor/sha_core/n3861_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_123 ),
	.I3(\top/processor/sha_core/n3489_159 ),
	.F(\top/processor/sha_core/n3861_107 )
);
defparam \top/processor/sha_core/n3861_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s180  (
	.I0(\top/processor/sha_core/n3503_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_149 ),
	.I3(\top/processor/sha_core/n3503_150 ),
	.F(\top/processor/sha_core/n3503_133 )
);
defparam \top/processor/sha_core/n3503_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s132  (
	.I0(\top/processor/sha_core/n3875_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_117 ),
	.I3(\top/processor/sha_core/n3503_150 ),
	.F(\top/processor/sha_core/n3875_101 )
);
defparam \top/processor/sha_core/n3875_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s181  (
	.I0(\top/processor/sha_core/n3503_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_152 ),
	.I3(\top/processor/sha_core/n3503_153 ),
	.F(\top/processor/sha_core/n3503_135 )
);
defparam \top/processor/sha_core/n3503_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s133  (
	.I0(\top/processor/sha_core/n3875_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_119 ),
	.I3(\top/processor/sha_core/n3503_153 ),
	.F(\top/processor/sha_core/n3875_103 )
);
defparam \top/processor/sha_core/n3875_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s182  (
	.I0(\top/processor/sha_core/n3503_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_155 ),
	.I3(\top/processor/sha_core/n3503_156 ),
	.F(\top/processor/sha_core/n3503_137 )
);
defparam \top/processor/sha_core/n3503_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s134  (
	.I0(\top/processor/sha_core/n3875_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_121 ),
	.I3(\top/processor/sha_core/n3503_156 ),
	.F(\top/processor/sha_core/n3875_105 )
);
defparam \top/processor/sha_core/n3875_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s183  (
	.I0(\top/processor/sha_core/n3503_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_158 ),
	.I3(\top/processor/sha_core/n3503_159 ),
	.F(\top/processor/sha_core/n3503_139 )
);
defparam \top/processor/sha_core/n3503_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s135  (
	.I0(\top/processor/sha_core/n3875_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_123 ),
	.I3(\top/processor/sha_core/n3503_159 ),
	.F(\top/processor/sha_core/n3875_107 )
);
defparam \top/processor/sha_core/n3875_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s184  (
	.I0(\top/processor/sha_core/n3503_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_161 ),
	.I3(\top/processor/sha_core/n3503_162 ),
	.F(\top/processor/sha_core/n3503_141 )
);
defparam \top/processor/sha_core/n3503_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s136  (
	.I0(\top/processor/sha_core/n3875_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_125 ),
	.I3(\top/processor/sha_core/n3503_162 ),
	.F(\top/processor/sha_core/n3875_109 )
);
defparam \top/processor/sha_core/n3875_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s185  (
	.I0(\top/processor/sha_core/n3503_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_164 ),
	.I3(\top/processor/sha_core/n3503_165 ),
	.F(\top/processor/sha_core/n3503_143 )
);
defparam \top/processor/sha_core/n3503_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s137  (
	.I0(\top/processor/sha_core/n3875_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_127 ),
	.I3(\top/processor/sha_core/n3503_165 ),
	.F(\top/processor/sha_core/n3875_111 )
);
defparam \top/processor/sha_core/n3875_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s186  (
	.I0(\top/processor/sha_core/n3503_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_167 ),
	.I3(\top/processor/sha_core/n3503_168 ),
	.F(\top/processor/sha_core/n3503_145 )
);
defparam \top/processor/sha_core/n3503_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s138  (
	.I0(\top/processor/sha_core/n3875_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_129 ),
	.I3(\top/processor/sha_core/n3503_168 ),
	.F(\top/processor/sha_core/n3875_113 )
);
defparam \top/processor/sha_core/n3875_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3503_s187  (
	.I0(\top/processor/sha_core/n3503_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_170 ),
	.I3(\top/processor/sha_core/n3503_171 ),
	.F(\top/processor/sha_core/n3503_147 )
);
defparam \top/processor/sha_core/n3503_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3875_s139  (
	.I0(\top/processor/sha_core/n3875_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3875_131 ),
	.I3(\top/processor/sha_core/n3503_171 ),
	.F(\top/processor/sha_core/n3875_115 )
);
defparam \top/processor/sha_core/n3875_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s180  (
	.I0(\top/processor/sha_core/n3504_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_149 ),
	.I3(\top/processor/sha_core/n3504_150 ),
	.F(\top/processor/sha_core/n3504_133 )
);
defparam \top/processor/sha_core/n3504_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s132  (
	.I0(\top/processor/sha_core/n3876_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_117 ),
	.I3(\top/processor/sha_core/n3504_150 ),
	.F(\top/processor/sha_core/n3876_101 )
);
defparam \top/processor/sha_core/n3876_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s181  (
	.I0(\top/processor/sha_core/n3504_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_152 ),
	.I3(\top/processor/sha_core/n3504_153 ),
	.F(\top/processor/sha_core/n3504_135 )
);
defparam \top/processor/sha_core/n3504_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s133  (
	.I0(\top/processor/sha_core/n3876_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_119 ),
	.I3(\top/processor/sha_core/n3504_153 ),
	.F(\top/processor/sha_core/n3876_103 )
);
defparam \top/processor/sha_core/n3876_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s184  (
	.I0(\top/processor/sha_core/n3489_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_161 ),
	.I3(\top/processor/sha_core/n3489_162 ),
	.F(\top/processor/sha_core/n3489_141 )
);
defparam \top/processor/sha_core/n3489_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s136  (
	.I0(\top/processor/sha_core/n3861_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_125 ),
	.I3(\top/processor/sha_core/n3489_162 ),
	.F(\top/processor/sha_core/n3861_109 )
);
defparam \top/processor/sha_core/n3861_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s182  (
	.I0(\top/processor/sha_core/n3504_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_155 ),
	.I3(\top/processor/sha_core/n3504_156 ),
	.F(\top/processor/sha_core/n3504_137 )
);
defparam \top/processor/sha_core/n3504_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s134  (
	.I0(\top/processor/sha_core/n3876_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_121 ),
	.I3(\top/processor/sha_core/n3504_156 ),
	.F(\top/processor/sha_core/n3876_105 )
);
defparam \top/processor/sha_core/n3876_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s183  (
	.I0(\top/processor/sha_core/n3504_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_158 ),
	.I3(\top/processor/sha_core/n3504_159 ),
	.F(\top/processor/sha_core/n3504_139 )
);
defparam \top/processor/sha_core/n3504_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s135  (
	.I0(\top/processor/sha_core/n3876_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_123 ),
	.I3(\top/processor/sha_core/n3504_159 ),
	.F(\top/processor/sha_core/n3876_107 )
);
defparam \top/processor/sha_core/n3876_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s184  (
	.I0(\top/processor/sha_core/n3504_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_161 ),
	.I3(\top/processor/sha_core/n3504_162 ),
	.F(\top/processor/sha_core/n3504_141 )
);
defparam \top/processor/sha_core/n3504_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s136  (
	.I0(\top/processor/sha_core/n3876_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_125 ),
	.I3(\top/processor/sha_core/n3504_162 ),
	.F(\top/processor/sha_core/n3876_109 )
);
defparam \top/processor/sha_core/n3876_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s185  (
	.I0(\top/processor/sha_core/n3504_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_164 ),
	.I3(\top/processor/sha_core/n3504_165 ),
	.F(\top/processor/sha_core/n3504_143 )
);
defparam \top/processor/sha_core/n3504_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s137  (
	.I0(\top/processor/sha_core/n3876_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_127 ),
	.I3(\top/processor/sha_core/n3504_165 ),
	.F(\top/processor/sha_core/n3876_111 )
);
defparam \top/processor/sha_core/n3876_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s186  (
	.I0(\top/processor/sha_core/n3504_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_167 ),
	.I3(\top/processor/sha_core/n3504_168 ),
	.F(\top/processor/sha_core/n3504_145 )
);
defparam \top/processor/sha_core/n3504_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s138  (
	.I0(\top/processor/sha_core/n3876_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_129 ),
	.I3(\top/processor/sha_core/n3504_168 ),
	.F(\top/processor/sha_core/n3876_113 )
);
defparam \top/processor/sha_core/n3876_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3504_s187  (
	.I0(\top/processor/sha_core/n3504_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_170 ),
	.I3(\top/processor/sha_core/n3504_171 ),
	.F(\top/processor/sha_core/n3504_147 )
);
defparam \top/processor/sha_core/n3504_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3876_s139  (
	.I0(\top/processor/sha_core/n3876_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3876_131 ),
	.I3(\top/processor/sha_core/n3504_171 ),
	.F(\top/processor/sha_core/n3876_115 )
);
defparam \top/processor/sha_core/n3876_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s180  (
	.I0(\top/processor/sha_core/n3505_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_149 ),
	.I3(\top/processor/sha_core/n3505_150 ),
	.F(\top/processor/sha_core/n3505_133 )
);
defparam \top/processor/sha_core/n3505_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s132  (
	.I0(\top/processor/sha_core/n3877_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_117 ),
	.I3(\top/processor/sha_core/n3505_150 ),
	.F(\top/processor/sha_core/n3877_101 )
);
defparam \top/processor/sha_core/n3877_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s181  (
	.I0(\top/processor/sha_core/n3505_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_152 ),
	.I3(\top/processor/sha_core/n3505_153 ),
	.F(\top/processor/sha_core/n3505_135 )
);
defparam \top/processor/sha_core/n3505_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s133  (
	.I0(\top/processor/sha_core/n3877_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_119 ),
	.I3(\top/processor/sha_core/n3505_153 ),
	.F(\top/processor/sha_core/n3877_103 )
);
defparam \top/processor/sha_core/n3877_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s182  (
	.I0(\top/processor/sha_core/n3505_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_155 ),
	.I3(\top/processor/sha_core/n3505_156 ),
	.F(\top/processor/sha_core/n3505_137 )
);
defparam \top/processor/sha_core/n3505_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s134  (
	.I0(\top/processor/sha_core/n3877_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_121 ),
	.I3(\top/processor/sha_core/n3505_156 ),
	.F(\top/processor/sha_core/n3877_105 )
);
defparam \top/processor/sha_core/n3877_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s183  (
	.I0(\top/processor/sha_core/n3505_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_158 ),
	.I3(\top/processor/sha_core/n3505_159 ),
	.F(\top/processor/sha_core/n3505_139 )
);
defparam \top/processor/sha_core/n3505_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s135  (
	.I0(\top/processor/sha_core/n3877_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_123 ),
	.I3(\top/processor/sha_core/n3505_159 ),
	.F(\top/processor/sha_core/n3877_107 )
);
defparam \top/processor/sha_core/n3877_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s185  (
	.I0(\top/processor/sha_core/n3489_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_164 ),
	.I3(\top/processor/sha_core/n3489_165 ),
	.F(\top/processor/sha_core/n3489_143 )
);
defparam \top/processor/sha_core/n3489_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s137  (
	.I0(\top/processor/sha_core/n3861_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_127 ),
	.I3(\top/processor/sha_core/n3489_165 ),
	.F(\top/processor/sha_core/n3861_111 )
);
defparam \top/processor/sha_core/n3861_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s184  (
	.I0(\top/processor/sha_core/n3505_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_161 ),
	.I3(\top/processor/sha_core/n3505_162 ),
	.F(\top/processor/sha_core/n3505_141 )
);
defparam \top/processor/sha_core/n3505_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s136  (
	.I0(\top/processor/sha_core/n3877_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_125 ),
	.I3(\top/processor/sha_core/n3505_162 ),
	.F(\top/processor/sha_core/n3877_109 )
);
defparam \top/processor/sha_core/n3877_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s185  (
	.I0(\top/processor/sha_core/n3505_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_164 ),
	.I3(\top/processor/sha_core/n3505_165 ),
	.F(\top/processor/sha_core/n3505_143 )
);
defparam \top/processor/sha_core/n3505_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s137  (
	.I0(\top/processor/sha_core/n3877_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_127 ),
	.I3(\top/processor/sha_core/n3505_165 ),
	.F(\top/processor/sha_core/n3877_111 )
);
defparam \top/processor/sha_core/n3877_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s186  (
	.I0(\top/processor/sha_core/n3505_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_167 ),
	.I3(\top/processor/sha_core/n3505_168 ),
	.F(\top/processor/sha_core/n3505_145 )
);
defparam \top/processor/sha_core/n3505_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s138  (
	.I0(\top/processor/sha_core/n3877_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_129 ),
	.I3(\top/processor/sha_core/n3505_168 ),
	.F(\top/processor/sha_core/n3877_113 )
);
defparam \top/processor/sha_core/n3877_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3505_s187  (
	.I0(\top/processor/sha_core/n3505_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_170 ),
	.I3(\top/processor/sha_core/n3505_171 ),
	.F(\top/processor/sha_core/n3505_147 )
);
defparam \top/processor/sha_core/n3505_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3877_s139  (
	.I0(\top/processor/sha_core/n3877_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3877_131 ),
	.I3(\top/processor/sha_core/n3505_171 ),
	.F(\top/processor/sha_core/n3877_115 )
);
defparam \top/processor/sha_core/n3877_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s180  (
	.I0(\top/processor/sha_core/n3506_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_149 ),
	.I3(\top/processor/sha_core/n3506_150 ),
	.F(\top/processor/sha_core/n3506_133 )
);
defparam \top/processor/sha_core/n3506_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s132  (
	.I0(\top/processor/sha_core/n3878_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_117 ),
	.I3(\top/processor/sha_core/n3506_150 ),
	.F(\top/processor/sha_core/n3878_101 )
);
defparam \top/processor/sha_core/n3878_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s181  (
	.I0(\top/processor/sha_core/n3506_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_152 ),
	.I3(\top/processor/sha_core/n3506_153 ),
	.F(\top/processor/sha_core/n3506_135 )
);
defparam \top/processor/sha_core/n3506_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s133  (
	.I0(\top/processor/sha_core/n3878_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_119 ),
	.I3(\top/processor/sha_core/n3506_153 ),
	.F(\top/processor/sha_core/n3878_103 )
);
defparam \top/processor/sha_core/n3878_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s182  (
	.I0(\top/processor/sha_core/n3506_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_155 ),
	.I3(\top/processor/sha_core/n3506_156 ),
	.F(\top/processor/sha_core/n3506_137 )
);
defparam \top/processor/sha_core/n3506_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s134  (
	.I0(\top/processor/sha_core/n3878_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_121 ),
	.I3(\top/processor/sha_core/n3506_156 ),
	.F(\top/processor/sha_core/n3878_105 )
);
defparam \top/processor/sha_core/n3878_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s183  (
	.I0(\top/processor/sha_core/n3506_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_158 ),
	.I3(\top/processor/sha_core/n3506_159 ),
	.F(\top/processor/sha_core/n3506_139 )
);
defparam \top/processor/sha_core/n3506_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s135  (
	.I0(\top/processor/sha_core/n3878_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_123 ),
	.I3(\top/processor/sha_core/n3506_159 ),
	.F(\top/processor/sha_core/n3878_107 )
);
defparam \top/processor/sha_core/n3878_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s184  (
	.I0(\top/processor/sha_core/n3506_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_161 ),
	.I3(\top/processor/sha_core/n3506_162 ),
	.F(\top/processor/sha_core/n3506_141 )
);
defparam \top/processor/sha_core/n3506_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s136  (
	.I0(\top/processor/sha_core/n3878_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_125 ),
	.I3(\top/processor/sha_core/n3506_162 ),
	.F(\top/processor/sha_core/n3878_109 )
);
defparam \top/processor/sha_core/n3878_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s185  (
	.I0(\top/processor/sha_core/n3506_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_164 ),
	.I3(\top/processor/sha_core/n3506_165 ),
	.F(\top/processor/sha_core/n3506_143 )
);
defparam \top/processor/sha_core/n3506_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s137  (
	.I0(\top/processor/sha_core/n3878_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_127 ),
	.I3(\top/processor/sha_core/n3506_165 ),
	.F(\top/processor/sha_core/n3878_111 )
);
defparam \top/processor/sha_core/n3878_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s186  (
	.I0(\top/processor/sha_core/n3489_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_167 ),
	.I3(\top/processor/sha_core/n3489_168 ),
	.F(\top/processor/sha_core/n3489_145 )
);
defparam \top/processor/sha_core/n3489_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s138  (
	.I0(\top/processor/sha_core/n3861_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_129 ),
	.I3(\top/processor/sha_core/n3489_168 ),
	.F(\top/processor/sha_core/n3861_113 )
);
defparam \top/processor/sha_core/n3861_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s186  (
	.I0(\top/processor/sha_core/n3506_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_167 ),
	.I3(\top/processor/sha_core/n3506_168 ),
	.F(\top/processor/sha_core/n3506_145 )
);
defparam \top/processor/sha_core/n3506_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s138  (
	.I0(\top/processor/sha_core/n3878_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_129 ),
	.I3(\top/processor/sha_core/n3506_168 ),
	.F(\top/processor/sha_core/n3878_113 )
);
defparam \top/processor/sha_core/n3878_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3506_s187  (
	.I0(\top/processor/sha_core/n3506_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_170 ),
	.I3(\top/processor/sha_core/n3506_171 ),
	.F(\top/processor/sha_core/n3506_147 )
);
defparam \top/processor/sha_core/n3506_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3878_s139  (
	.I0(\top/processor/sha_core/n3878_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3878_131 ),
	.I3(\top/processor/sha_core/n3506_171 ),
	.F(\top/processor/sha_core/n3878_115 )
);
defparam \top/processor/sha_core/n3878_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s180  (
	.I0(\top/processor/sha_core/n3507_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_149 ),
	.I3(\top/processor/sha_core/n3507_150 ),
	.F(\top/processor/sha_core/n3507_133 )
);
defparam \top/processor/sha_core/n3507_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s132  (
	.I0(\top/processor/sha_core/n3879_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_117 ),
	.I3(\top/processor/sha_core/n3507_150 ),
	.F(\top/processor/sha_core/n3879_101 )
);
defparam \top/processor/sha_core/n3879_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s181  (
	.I0(\top/processor/sha_core/n3507_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_152 ),
	.I3(\top/processor/sha_core/n3507_153 ),
	.F(\top/processor/sha_core/n3507_135 )
);
defparam \top/processor/sha_core/n3507_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s133  (
	.I0(\top/processor/sha_core/n3879_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_119 ),
	.I3(\top/processor/sha_core/n3507_153 ),
	.F(\top/processor/sha_core/n3879_103 )
);
defparam \top/processor/sha_core/n3879_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s182  (
	.I0(\top/processor/sha_core/n3507_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_155 ),
	.I3(\top/processor/sha_core/n3507_156 ),
	.F(\top/processor/sha_core/n3507_137 )
);
defparam \top/processor/sha_core/n3507_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s134  (
	.I0(\top/processor/sha_core/n3879_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_121 ),
	.I3(\top/processor/sha_core/n3507_156 ),
	.F(\top/processor/sha_core/n3879_105 )
);
defparam \top/processor/sha_core/n3879_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s183  (
	.I0(\top/processor/sha_core/n3507_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_158 ),
	.I3(\top/processor/sha_core/n3507_159 ),
	.F(\top/processor/sha_core/n3507_139 )
);
defparam \top/processor/sha_core/n3507_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s135  (
	.I0(\top/processor/sha_core/n3879_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_123 ),
	.I3(\top/processor/sha_core/n3507_159 ),
	.F(\top/processor/sha_core/n3879_107 )
);
defparam \top/processor/sha_core/n3879_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s184  (
	.I0(\top/processor/sha_core/n3507_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_161 ),
	.I3(\top/processor/sha_core/n3507_162 ),
	.F(\top/processor/sha_core/n3507_141 )
);
defparam \top/processor/sha_core/n3507_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s136  (
	.I0(\top/processor/sha_core/n3879_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_125 ),
	.I3(\top/processor/sha_core/n3507_162 ),
	.F(\top/processor/sha_core/n3879_109 )
);
defparam \top/processor/sha_core/n3879_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s185  (
	.I0(\top/processor/sha_core/n3507_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_164 ),
	.I3(\top/processor/sha_core/n3507_165 ),
	.F(\top/processor/sha_core/n3507_143 )
);
defparam \top/processor/sha_core/n3507_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s137  (
	.I0(\top/processor/sha_core/n3879_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_127 ),
	.I3(\top/processor/sha_core/n3507_165 ),
	.F(\top/processor/sha_core/n3879_111 )
);
defparam \top/processor/sha_core/n3879_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s186  (
	.I0(\top/processor/sha_core/n3507_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_167 ),
	.I3(\top/processor/sha_core/n3507_168 ),
	.F(\top/processor/sha_core/n3507_145 )
);
defparam \top/processor/sha_core/n3507_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s138  (
	.I0(\top/processor/sha_core/n3879_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_129 ),
	.I3(\top/processor/sha_core/n3507_168 ),
	.F(\top/processor/sha_core/n3879_113 )
);
defparam \top/processor/sha_core/n3879_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3507_s187  (
	.I0(\top/processor/sha_core/n3507_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_170 ),
	.I3(\top/processor/sha_core/n3507_171 ),
	.F(\top/processor/sha_core/n3507_147 )
);
defparam \top/processor/sha_core/n3507_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3879_s139  (
	.I0(\top/processor/sha_core/n3879_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3879_131 ),
	.I3(\top/processor/sha_core/n3507_171 ),
	.F(\top/processor/sha_core/n3879_115 )
);
defparam \top/processor/sha_core/n3879_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3489_s187  (
	.I0(\top/processor/sha_core/n3489_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_170 ),
	.I3(\top/processor/sha_core/n3489_171 ),
	.F(\top/processor/sha_core/n3489_147 )
);
defparam \top/processor/sha_core/n3489_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3861_s139  (
	.I0(\top/processor/sha_core/n3861_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3861_131 ),
	.I3(\top/processor/sha_core/n3489_171 ),
	.F(\top/processor/sha_core/n3861_115 )
);
defparam \top/processor/sha_core/n3861_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s180  (
	.I0(\top/processor/sha_core/n3508_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_149 ),
	.I3(\top/processor/sha_core/n3508_150 ),
	.F(\top/processor/sha_core/n3508_133 )
);
defparam \top/processor/sha_core/n3508_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s132  (
	.I0(\top/processor/sha_core/n3880_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_117 ),
	.I3(\top/processor/sha_core/n3508_150 ),
	.F(\top/processor/sha_core/n3880_101 )
);
defparam \top/processor/sha_core/n3880_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s181  (
	.I0(\top/processor/sha_core/n3508_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_152 ),
	.I3(\top/processor/sha_core/n3508_153 ),
	.F(\top/processor/sha_core/n3508_135 )
);
defparam \top/processor/sha_core/n3508_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s133  (
	.I0(\top/processor/sha_core/n3880_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_119 ),
	.I3(\top/processor/sha_core/n3508_153 ),
	.F(\top/processor/sha_core/n3880_103 )
);
defparam \top/processor/sha_core/n3880_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s182  (
	.I0(\top/processor/sha_core/n3508_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_155 ),
	.I3(\top/processor/sha_core/n3508_156 ),
	.F(\top/processor/sha_core/n3508_137 )
);
defparam \top/processor/sha_core/n3508_s182 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3880_s134  (
	.I0(\top/processor/sha_core/n3880_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_121 ),
	.I3(\top/processor/sha_core/n3508_156 ),
	.F(\top/processor/sha_core/n3880_105 )
);
defparam \top/processor/sha_core/n3880_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s183  (
	.I0(\top/processor/sha_core/n3508_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_158 ),
	.I3(\top/processor/sha_core/n3508_159 ),
	.F(\top/processor/sha_core/n3508_139 )
);
defparam \top/processor/sha_core/n3508_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s135  (
	.I0(\top/processor/sha_core/n3880_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_123 ),
	.I3(\top/processor/sha_core/n3508_159 ),
	.F(\top/processor/sha_core/n3880_107 )
);
defparam \top/processor/sha_core/n3880_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s184  (
	.I0(\top/processor/sha_core/n3508_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_161 ),
	.I3(\top/processor/sha_core/n3508_162 ),
	.F(\top/processor/sha_core/n3508_141 )
);
defparam \top/processor/sha_core/n3508_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s136  (
	.I0(\top/processor/sha_core/n3880_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_125 ),
	.I3(\top/processor/sha_core/n3508_162 ),
	.F(\top/processor/sha_core/n3880_109 )
);
defparam \top/processor/sha_core/n3880_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s185  (
	.I0(\top/processor/sha_core/n3508_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_164 ),
	.I3(\top/processor/sha_core/n3508_165 ),
	.F(\top/processor/sha_core/n3508_143 )
);
defparam \top/processor/sha_core/n3508_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s137  (
	.I0(\top/processor/sha_core/n3880_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_127 ),
	.I3(\top/processor/sha_core/n3508_165 ),
	.F(\top/processor/sha_core/n3880_111 )
);
defparam \top/processor/sha_core/n3880_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s186  (
	.I0(\top/processor/sha_core/n3508_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_167 ),
	.I3(\top/processor/sha_core/n3508_168 ),
	.F(\top/processor/sha_core/n3508_145 )
);
defparam \top/processor/sha_core/n3508_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s138  (
	.I0(\top/processor/sha_core/n3880_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_129 ),
	.I3(\top/processor/sha_core/n3508_168 ),
	.F(\top/processor/sha_core/n3880_113 )
);
defparam \top/processor/sha_core/n3880_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3508_s187  (
	.I0(\top/processor/sha_core/n3508_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_170 ),
	.I3(\top/processor/sha_core/n3508_171 ),
	.F(\top/processor/sha_core/n3508_147 )
);
defparam \top/processor/sha_core/n3508_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3880_s139  (
	.I0(\top/processor/sha_core/n3880_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3880_131 ),
	.I3(\top/processor/sha_core/n3508_171 ),
	.F(\top/processor/sha_core/n3880_115 )
);
defparam \top/processor/sha_core/n3880_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3509_s180  (
	.I0(\top/processor/sha_core/n3509_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_149 ),
	.I3(\top/processor/sha_core/n3509_150 ),
	.F(\top/processor/sha_core/n3509_133 )
);
defparam \top/processor/sha_core/n3509_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s132  (
	.I0(\top/processor/sha_core/n3881_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_117 ),
	.I3(\top/processor/sha_core/n3509_150 ),
	.F(\top/processor/sha_core/n3881_101 )
);
defparam \top/processor/sha_core/n3881_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s181  (
	.I0(\top/processor/sha_core/n3509_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_152 ),
	.I3(\top/processor/sha_core/n3509_153 ),
	.F(\top/processor/sha_core/n3509_135 )
);
defparam \top/processor/sha_core/n3509_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s133  (
	.I0(\top/processor/sha_core/n3881_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_119 ),
	.I3(\top/processor/sha_core/n3509_153 ),
	.F(\top/processor/sha_core/n3881_103 )
);
defparam \top/processor/sha_core/n3881_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s180  (
	.I0(\top/processor/sha_core/n3490_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_149 ),
	.I3(\top/processor/sha_core/n3490_150 ),
	.F(\top/processor/sha_core/n3490_133 )
);
defparam \top/processor/sha_core/n3490_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s132  (
	.I0(\top/processor/sha_core/n3862_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_117 ),
	.I3(\top/processor/sha_core/n3490_150 ),
	.F(\top/processor/sha_core/n3862_101 )
);
defparam \top/processor/sha_core/n3862_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s182  (
	.I0(\top/processor/sha_core/n3509_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_155 ),
	.I3(\top/processor/sha_core/n3509_156 ),
	.F(\top/processor/sha_core/n3509_137 )
);
defparam \top/processor/sha_core/n3509_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s134  (
	.I0(\top/processor/sha_core/n3881_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_121 ),
	.I3(\top/processor/sha_core/n3509_156 ),
	.F(\top/processor/sha_core/n3881_105 )
);
defparam \top/processor/sha_core/n3881_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s183  (
	.I0(\top/processor/sha_core/n3509_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_158 ),
	.I3(\top/processor/sha_core/n3509_159 ),
	.F(\top/processor/sha_core/n3509_139 )
);
defparam \top/processor/sha_core/n3509_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s135  (
	.I0(\top/processor/sha_core/n3881_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_123 ),
	.I3(\top/processor/sha_core/n3509_159 ),
	.F(\top/processor/sha_core/n3881_107 )
);
defparam \top/processor/sha_core/n3881_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s184  (
	.I0(\top/processor/sha_core/n3509_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_161 ),
	.I3(\top/processor/sha_core/n3509_162 ),
	.F(\top/processor/sha_core/n3509_141 )
);
defparam \top/processor/sha_core/n3509_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s136  (
	.I0(\top/processor/sha_core/n3881_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_125 ),
	.I3(\top/processor/sha_core/n3509_162 ),
	.F(\top/processor/sha_core/n3881_109 )
);
defparam \top/processor/sha_core/n3881_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s185  (
	.I0(\top/processor/sha_core/n3509_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_164 ),
	.I3(\top/processor/sha_core/n3509_165 ),
	.F(\top/processor/sha_core/n3509_143 )
);
defparam \top/processor/sha_core/n3509_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s137  (
	.I0(\top/processor/sha_core/n3881_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_127 ),
	.I3(\top/processor/sha_core/n3509_165 ),
	.F(\top/processor/sha_core/n3881_111 )
);
defparam \top/processor/sha_core/n3881_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s186  (
	.I0(\top/processor/sha_core/n3509_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_167 ),
	.I3(\top/processor/sha_core/n3509_168 ),
	.F(\top/processor/sha_core/n3509_145 )
);
defparam \top/processor/sha_core/n3509_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s138  (
	.I0(\top/processor/sha_core/n3881_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_129 ),
	.I3(\top/processor/sha_core/n3509_168 ),
	.F(\top/processor/sha_core/n3881_113 )
);
defparam \top/processor/sha_core/n3881_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3509_s187  (
	.I0(\top/processor/sha_core/n3509_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_170 ),
	.I3(\top/processor/sha_core/n3509_171 ),
	.F(\top/processor/sha_core/n3509_147 )
);
defparam \top/processor/sha_core/n3509_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3881_s139  (
	.I0(\top/processor/sha_core/n3881_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3881_131 ),
	.I3(\top/processor/sha_core/n3509_171 ),
	.F(\top/processor/sha_core/n3881_115 )
);
defparam \top/processor/sha_core/n3881_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s180  (
	.I0(\top/processor/sha_core/n3510_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_149 ),
	.I3(\top/processor/sha_core/n3510_150 ),
	.F(\top/processor/sha_core/n3510_133 )
);
defparam \top/processor/sha_core/n3510_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s132  (
	.I0(\top/processor/sha_core/n3882_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_117 ),
	.I3(\top/processor/sha_core/n3510_150 ),
	.F(\top/processor/sha_core/n3882_101 )
);
defparam \top/processor/sha_core/n3882_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s181  (
	.I0(\top/processor/sha_core/n3510_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_152 ),
	.I3(\top/processor/sha_core/n3510_153 ),
	.F(\top/processor/sha_core/n3510_135 )
);
defparam \top/processor/sha_core/n3510_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s133  (
	.I0(\top/processor/sha_core/n3882_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_119 ),
	.I3(\top/processor/sha_core/n3510_153 ),
	.F(\top/processor/sha_core/n3882_103 )
);
defparam \top/processor/sha_core/n3882_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s182  (
	.I0(\top/processor/sha_core/n3510_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_155 ),
	.I3(\top/processor/sha_core/n3510_156 ),
	.F(\top/processor/sha_core/n3510_137 )
);
defparam \top/processor/sha_core/n3510_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s134  (
	.I0(\top/processor/sha_core/n3882_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_121 ),
	.I3(\top/processor/sha_core/n3510_156 ),
	.F(\top/processor/sha_core/n3882_105 )
);
defparam \top/processor/sha_core/n3882_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s183  (
	.I0(\top/processor/sha_core/n3510_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_158 ),
	.I3(\top/processor/sha_core/n3510_159 ),
	.F(\top/processor/sha_core/n3510_139 )
);
defparam \top/processor/sha_core/n3510_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s135  (
	.I0(\top/processor/sha_core/n3882_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_123 ),
	.I3(\top/processor/sha_core/n3510_159 ),
	.F(\top/processor/sha_core/n3882_107 )
);
defparam \top/processor/sha_core/n3882_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s181  (
	.I0(\top/processor/sha_core/n3490_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_152 ),
	.I3(\top/processor/sha_core/n3490_153 ),
	.F(\top/processor/sha_core/n3490_135 )
);
defparam \top/processor/sha_core/n3490_s181 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3862_s133  (
	.I0(\top/processor/sha_core/n3862_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_119 ),
	.I3(\top/processor/sha_core/n3490_153 ),
	.F(\top/processor/sha_core/n3862_103 )
);
defparam \top/processor/sha_core/n3862_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s184  (
	.I0(\top/processor/sha_core/n3510_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_161 ),
	.I3(\top/processor/sha_core/n3510_162 ),
	.F(\top/processor/sha_core/n3510_141 )
);
defparam \top/processor/sha_core/n3510_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s136  (
	.I0(\top/processor/sha_core/n3882_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_125 ),
	.I3(\top/processor/sha_core/n3510_162 ),
	.F(\top/processor/sha_core/n3882_109 )
);
defparam \top/processor/sha_core/n3882_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s185  (
	.I0(\top/processor/sha_core/n3510_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_164 ),
	.I3(\top/processor/sha_core/n3510_165 ),
	.F(\top/processor/sha_core/n3510_143 )
);
defparam \top/processor/sha_core/n3510_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s137  (
	.I0(\top/processor/sha_core/n3882_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_127 ),
	.I3(\top/processor/sha_core/n3510_165 ),
	.F(\top/processor/sha_core/n3882_111 )
);
defparam \top/processor/sha_core/n3882_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s186  (
	.I0(\top/processor/sha_core/n3510_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_167 ),
	.I3(\top/processor/sha_core/n3510_168 ),
	.F(\top/processor/sha_core/n3510_145 )
);
defparam \top/processor/sha_core/n3510_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s138  (
	.I0(\top/processor/sha_core/n3882_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_129 ),
	.I3(\top/processor/sha_core/n3510_168 ),
	.F(\top/processor/sha_core/n3882_113 )
);
defparam \top/processor/sha_core/n3882_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3510_s187  (
	.I0(\top/processor/sha_core/n3510_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_170 ),
	.I3(\top/processor/sha_core/n3510_171 ),
	.F(\top/processor/sha_core/n3510_147 )
);
defparam \top/processor/sha_core/n3510_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3882_s139  (
	.I0(\top/processor/sha_core/n3882_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3882_131 ),
	.I3(\top/processor/sha_core/n3510_171 ),
	.F(\top/processor/sha_core/n3882_115 )
);
defparam \top/processor/sha_core/n3882_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s180  (
	.I0(\top/processor/sha_core/n3511_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_149 ),
	.I3(\top/processor/sha_core/n3511_150 ),
	.F(\top/processor/sha_core/n3511_133 )
);
defparam \top/processor/sha_core/n3511_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s132  (
	.I0(\top/processor/sha_core/n3883_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_117 ),
	.I3(\top/processor/sha_core/n3511_150 ),
	.F(\top/processor/sha_core/n3883_101 )
);
defparam \top/processor/sha_core/n3883_s132 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3511_s181  (
	.I0(\top/processor/sha_core/n3511_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_152 ),
	.I3(\top/processor/sha_core/n3511_153 ),
	.F(\top/processor/sha_core/n3511_135 )
);
defparam \top/processor/sha_core/n3511_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s133  (
	.I0(\top/processor/sha_core/n3883_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_119 ),
	.I3(\top/processor/sha_core/n3511_153 ),
	.F(\top/processor/sha_core/n3883_103 )
);
defparam \top/processor/sha_core/n3883_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s182  (
	.I0(\top/processor/sha_core/n3511_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_155 ),
	.I3(\top/processor/sha_core/n3511_156 ),
	.F(\top/processor/sha_core/n3511_137 )
);
defparam \top/processor/sha_core/n3511_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s134  (
	.I0(\top/processor/sha_core/n3883_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_121 ),
	.I3(\top/processor/sha_core/n3511_156 ),
	.F(\top/processor/sha_core/n3883_105 )
);
defparam \top/processor/sha_core/n3883_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s183  (
	.I0(\top/processor/sha_core/n3511_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_158 ),
	.I3(\top/processor/sha_core/n3511_159 ),
	.F(\top/processor/sha_core/n3511_139 )
);
defparam \top/processor/sha_core/n3511_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s135  (
	.I0(\top/processor/sha_core/n3883_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_123 ),
	.I3(\top/processor/sha_core/n3511_159 ),
	.F(\top/processor/sha_core/n3883_107 )
);
defparam \top/processor/sha_core/n3883_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s184  (
	.I0(\top/processor/sha_core/n3511_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_161 ),
	.I3(\top/processor/sha_core/n3511_162 ),
	.F(\top/processor/sha_core/n3511_141 )
);
defparam \top/processor/sha_core/n3511_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s136  (
	.I0(\top/processor/sha_core/n3883_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_125 ),
	.I3(\top/processor/sha_core/n3511_162 ),
	.F(\top/processor/sha_core/n3883_109 )
);
defparam \top/processor/sha_core/n3883_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s185  (
	.I0(\top/processor/sha_core/n3511_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_164 ),
	.I3(\top/processor/sha_core/n3511_165 ),
	.F(\top/processor/sha_core/n3511_143 )
);
defparam \top/processor/sha_core/n3511_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s137  (
	.I0(\top/processor/sha_core/n3883_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_127 ),
	.I3(\top/processor/sha_core/n3511_165 ),
	.F(\top/processor/sha_core/n3883_111 )
);
defparam \top/processor/sha_core/n3883_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s182  (
	.I0(\top/processor/sha_core/n3490_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_155 ),
	.I3(\top/processor/sha_core/n3490_156 ),
	.F(\top/processor/sha_core/n3490_137 )
);
defparam \top/processor/sha_core/n3490_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s134  (
	.I0(\top/processor/sha_core/n3862_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_121 ),
	.I3(\top/processor/sha_core/n3490_156 ),
	.F(\top/processor/sha_core/n3862_105 )
);
defparam \top/processor/sha_core/n3862_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s186  (
	.I0(\top/processor/sha_core/n3511_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_167 ),
	.I3(\top/processor/sha_core/n3511_168 ),
	.F(\top/processor/sha_core/n3511_145 )
);
defparam \top/processor/sha_core/n3511_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s138  (
	.I0(\top/processor/sha_core/n3883_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_129 ),
	.I3(\top/processor/sha_core/n3511_168 ),
	.F(\top/processor/sha_core/n3883_113 )
);
defparam \top/processor/sha_core/n3883_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3511_s187  (
	.I0(\top/processor/sha_core/n3511_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_170 ),
	.I3(\top/processor/sha_core/n3511_171 ),
	.F(\top/processor/sha_core/n3511_147 )
);
defparam \top/processor/sha_core/n3511_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3883_s139  (
	.I0(\top/processor/sha_core/n3883_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3883_131 ),
	.I3(\top/processor/sha_core/n3511_171 ),
	.F(\top/processor/sha_core/n3883_115 )
);
defparam \top/processor/sha_core/n3883_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s180  (
	.I0(\top/processor/sha_core/n3512_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_149 ),
	.I3(\top/processor/sha_core/n3512_150 ),
	.F(\top/processor/sha_core/n3512_133 )
);
defparam \top/processor/sha_core/n3512_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s132  (
	.I0(\top/processor/sha_core/n3884_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_117 ),
	.I3(\top/processor/sha_core/n3512_150 ),
	.F(\top/processor/sha_core/n3884_101 )
);
defparam \top/processor/sha_core/n3884_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s181  (
	.I0(\top/processor/sha_core/n3512_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_152 ),
	.I3(\top/processor/sha_core/n3512_153 ),
	.F(\top/processor/sha_core/n3512_135 )
);
defparam \top/processor/sha_core/n3512_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s133  (
	.I0(\top/processor/sha_core/n3884_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_119 ),
	.I3(\top/processor/sha_core/n3512_153 ),
	.F(\top/processor/sha_core/n3884_103 )
);
defparam \top/processor/sha_core/n3884_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s182  (
	.I0(\top/processor/sha_core/n3512_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_155 ),
	.I3(\top/processor/sha_core/n3512_156 ),
	.F(\top/processor/sha_core/n3512_137 )
);
defparam \top/processor/sha_core/n3512_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s134  (
	.I0(\top/processor/sha_core/n3884_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_121 ),
	.I3(\top/processor/sha_core/n3512_156 ),
	.F(\top/processor/sha_core/n3884_105 )
);
defparam \top/processor/sha_core/n3884_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s183  (
	.I0(\top/processor/sha_core/n3512_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_158 ),
	.I3(\top/processor/sha_core/n3512_159 ),
	.F(\top/processor/sha_core/n3512_139 )
);
defparam \top/processor/sha_core/n3512_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s135  (
	.I0(\top/processor/sha_core/n3884_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_123 ),
	.I3(\top/processor/sha_core/n3512_159 ),
	.F(\top/processor/sha_core/n3884_107 )
);
defparam \top/processor/sha_core/n3884_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s184  (
	.I0(\top/processor/sha_core/n3512_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_161 ),
	.I3(\top/processor/sha_core/n3512_162 ),
	.F(\top/processor/sha_core/n3512_141 )
);
defparam \top/processor/sha_core/n3512_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s136  (
	.I0(\top/processor/sha_core/n3884_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_125 ),
	.I3(\top/processor/sha_core/n3512_162 ),
	.F(\top/processor/sha_core/n3884_109 )
);
defparam \top/processor/sha_core/n3884_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s185  (
	.I0(\top/processor/sha_core/n3512_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_164 ),
	.I3(\top/processor/sha_core/n3512_165 ),
	.F(\top/processor/sha_core/n3512_143 )
);
defparam \top/processor/sha_core/n3512_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s137  (
	.I0(\top/processor/sha_core/n3884_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_127 ),
	.I3(\top/processor/sha_core/n3512_165 ),
	.F(\top/processor/sha_core/n3884_111 )
);
defparam \top/processor/sha_core/n3884_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s186  (
	.I0(\top/processor/sha_core/n3512_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_167 ),
	.I3(\top/processor/sha_core/n3512_168 ),
	.F(\top/processor/sha_core/n3512_145 )
);
defparam \top/processor/sha_core/n3512_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s138  (
	.I0(\top/processor/sha_core/n3884_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_129 ),
	.I3(\top/processor/sha_core/n3512_168 ),
	.F(\top/processor/sha_core/n3884_113 )
);
defparam \top/processor/sha_core/n3884_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3512_s187  (
	.I0(\top/processor/sha_core/n3512_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_170 ),
	.I3(\top/processor/sha_core/n3512_171 ),
	.F(\top/processor/sha_core/n3512_147 )
);
defparam \top/processor/sha_core/n3512_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3884_s139  (
	.I0(\top/processor/sha_core/n3884_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3884_131 ),
	.I3(\top/processor/sha_core/n3512_171 ),
	.F(\top/processor/sha_core/n3884_115 )
);
defparam \top/processor/sha_core/n3884_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s183  (
	.I0(\top/processor/sha_core/n3490_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_158 ),
	.I3(\top/processor/sha_core/n3490_159 ),
	.F(\top/processor/sha_core/n3490_139 )
);
defparam \top/processor/sha_core/n3490_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s135  (
	.I0(\top/processor/sha_core/n3862_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_123 ),
	.I3(\top/processor/sha_core/n3490_159 ),
	.F(\top/processor/sha_core/n3862_107 )
);
defparam \top/processor/sha_core/n3862_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s181  (
	.I0(\top/processor/sha_core/n3488_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_161 ),
	.I3(\top/processor/sha_core/n3488_162 ),
	.F(\top/processor/sha_core/n3488_141 )
);
defparam \top/processor/sha_core/n3488_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s133  (
	.I0(\top/processor/sha_core/n3860_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_125 ),
	.I3(\top/processor/sha_core/n3488_162 ),
	.F(\top/processor/sha_core/n3860_109 )
);
defparam \top/processor/sha_core/n3860_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s180  (
	.I0(\top/processor/sha_core/n3513_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_149 ),
	.I3(\top/processor/sha_core/n3513_150 ),
	.F(\top/processor/sha_core/n3513_133 )
);
defparam \top/processor/sha_core/n3513_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s132  (
	.I0(\top/processor/sha_core/n3885_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_117 ),
	.I3(\top/processor/sha_core/n3513_150 ),
	.F(\top/processor/sha_core/n3885_101 )
);
defparam \top/processor/sha_core/n3885_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s181  (
	.I0(\top/processor/sha_core/n3513_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_152 ),
	.I3(\top/processor/sha_core/n3513_153 ),
	.F(\top/processor/sha_core/n3513_135 )
);
defparam \top/processor/sha_core/n3513_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s133  (
	.I0(\top/processor/sha_core/n3885_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_119 ),
	.I3(\top/processor/sha_core/n3513_153 ),
	.F(\top/processor/sha_core/n3885_103 )
);
defparam \top/processor/sha_core/n3885_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s182  (
	.I0(\top/processor/sha_core/n3513_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_155 ),
	.I3(\top/processor/sha_core/n3513_156 ),
	.F(\top/processor/sha_core/n3513_137 )
);
defparam \top/processor/sha_core/n3513_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s134  (
	.I0(\top/processor/sha_core/n3885_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_121 ),
	.I3(\top/processor/sha_core/n3513_156 ),
	.F(\top/processor/sha_core/n3885_105 )
);
defparam \top/processor/sha_core/n3885_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s183  (
	.I0(\top/processor/sha_core/n3513_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_158 ),
	.I3(\top/processor/sha_core/n3513_159 ),
	.F(\top/processor/sha_core/n3513_139 )
);
defparam \top/processor/sha_core/n3513_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s135  (
	.I0(\top/processor/sha_core/n3885_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_123 ),
	.I3(\top/processor/sha_core/n3513_159 ),
	.F(\top/processor/sha_core/n3885_107 )
);
defparam \top/processor/sha_core/n3885_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s184  (
	.I0(\top/processor/sha_core/n3513_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_161 ),
	.I3(\top/processor/sha_core/n3513_162 ),
	.F(\top/processor/sha_core/n3513_141 )
);
defparam \top/processor/sha_core/n3513_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s136  (
	.I0(\top/processor/sha_core/n3885_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_125 ),
	.I3(\top/processor/sha_core/n3513_162 ),
	.F(\top/processor/sha_core/n3885_109 )
);
defparam \top/processor/sha_core/n3885_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s185  (
	.I0(\top/processor/sha_core/n3513_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_164 ),
	.I3(\top/processor/sha_core/n3513_165 ),
	.F(\top/processor/sha_core/n3513_143 )
);
defparam \top/processor/sha_core/n3513_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s137  (
	.I0(\top/processor/sha_core/n3885_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_127 ),
	.I3(\top/processor/sha_core/n3513_165 ),
	.F(\top/processor/sha_core/n3885_111 )
);
defparam \top/processor/sha_core/n3885_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s186  (
	.I0(\top/processor/sha_core/n3513_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_167 ),
	.I3(\top/processor/sha_core/n3513_168 ),
	.F(\top/processor/sha_core/n3513_145 )
);
defparam \top/processor/sha_core/n3513_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s138  (
	.I0(\top/processor/sha_core/n3885_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_129 ),
	.I3(\top/processor/sha_core/n3513_168 ),
	.F(\top/processor/sha_core/n3885_113 )
);
defparam \top/processor/sha_core/n3885_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3513_s187  (
	.I0(\top/processor/sha_core/n3513_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_170 ),
	.I3(\top/processor/sha_core/n3513_171 ),
	.F(\top/processor/sha_core/n3513_147 )
);
defparam \top/processor/sha_core/n3513_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3885_s139  (
	.I0(\top/processor/sha_core/n3885_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3885_131 ),
	.I3(\top/processor/sha_core/n3513_171 ),
	.F(\top/processor/sha_core/n3885_115 )
);
defparam \top/processor/sha_core/n3885_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s180  (
	.I0(\top/processor/sha_core/n3514_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_149 ),
	.I3(\top/processor/sha_core/n3514_150 ),
	.F(\top/processor/sha_core/n3514_133 )
);
defparam \top/processor/sha_core/n3514_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s132  (
	.I0(\top/processor/sha_core/n3886_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_117 ),
	.I3(\top/processor/sha_core/n3514_150 ),
	.F(\top/processor/sha_core/n3886_101 )
);
defparam \top/processor/sha_core/n3886_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s181  (
	.I0(\top/processor/sha_core/n3514_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_152 ),
	.I3(\top/processor/sha_core/n3514_153 ),
	.F(\top/processor/sha_core/n3514_135 )
);
defparam \top/processor/sha_core/n3514_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s133  (
	.I0(\top/processor/sha_core/n3886_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_119 ),
	.I3(\top/processor/sha_core/n3514_153 ),
	.F(\top/processor/sha_core/n3886_103 )
);
defparam \top/processor/sha_core/n3886_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s184  (
	.I0(\top/processor/sha_core/n3490_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_161 ),
	.I3(\top/processor/sha_core/n3490_162 ),
	.F(\top/processor/sha_core/n3490_141 )
);
defparam \top/processor/sha_core/n3490_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s136  (
	.I0(\top/processor/sha_core/n3862_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_125 ),
	.I3(\top/processor/sha_core/n3490_162 ),
	.F(\top/processor/sha_core/n3862_109 )
);
defparam \top/processor/sha_core/n3862_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s182  (
	.I0(\top/processor/sha_core/n3514_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_155 ),
	.I3(\top/processor/sha_core/n3514_156 ),
	.F(\top/processor/sha_core/n3514_137 )
);
defparam \top/processor/sha_core/n3514_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s134  (
	.I0(\top/processor/sha_core/n3886_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_121 ),
	.I3(\top/processor/sha_core/n3514_156 ),
	.F(\top/processor/sha_core/n3886_105 )
);
defparam \top/processor/sha_core/n3886_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s183  (
	.I0(\top/processor/sha_core/n3514_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_158 ),
	.I3(\top/processor/sha_core/n3514_159 ),
	.F(\top/processor/sha_core/n3514_139 )
);
defparam \top/processor/sha_core/n3514_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s135  (
	.I0(\top/processor/sha_core/n3886_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_123 ),
	.I3(\top/processor/sha_core/n3514_159 ),
	.F(\top/processor/sha_core/n3886_107 )
);
defparam \top/processor/sha_core/n3886_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s184  (
	.I0(\top/processor/sha_core/n3514_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_161 ),
	.I3(\top/processor/sha_core/n3514_162 ),
	.F(\top/processor/sha_core/n3514_141 )
);
defparam \top/processor/sha_core/n3514_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s136  (
	.I0(\top/processor/sha_core/n3886_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_125 ),
	.I3(\top/processor/sha_core/n3514_162 ),
	.F(\top/processor/sha_core/n3886_109 )
);
defparam \top/processor/sha_core/n3886_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s185  (
	.I0(\top/processor/sha_core/n3514_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_164 ),
	.I3(\top/processor/sha_core/n3514_165 ),
	.F(\top/processor/sha_core/n3514_143 )
);
defparam \top/processor/sha_core/n3514_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s137  (
	.I0(\top/processor/sha_core/n3886_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_127 ),
	.I3(\top/processor/sha_core/n3514_165 ),
	.F(\top/processor/sha_core/n3886_111 )
);
defparam \top/processor/sha_core/n3886_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s186  (
	.I0(\top/processor/sha_core/n3514_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_167 ),
	.I3(\top/processor/sha_core/n3514_168 ),
	.F(\top/processor/sha_core/n3514_145 )
);
defparam \top/processor/sha_core/n3514_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s138  (
	.I0(\top/processor/sha_core/n3886_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_129 ),
	.I3(\top/processor/sha_core/n3514_168 ),
	.F(\top/processor/sha_core/n3886_113 )
);
defparam \top/processor/sha_core/n3886_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3514_s187  (
	.I0(\top/processor/sha_core/n3514_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_170 ),
	.I3(\top/processor/sha_core/n3514_171 ),
	.F(\top/processor/sha_core/n3514_147 )
);
defparam \top/processor/sha_core/n3514_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3886_s139  (
	.I0(\top/processor/sha_core/n3886_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3886_131 ),
	.I3(\top/processor/sha_core/n3514_171 ),
	.F(\top/processor/sha_core/n3886_115 )
);
defparam \top/processor/sha_core/n3886_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s180  (
	.I0(\top/processor/sha_core/n3515_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_149 ),
	.I3(\top/processor/sha_core/n3515_150 ),
	.F(\top/processor/sha_core/n3515_133 )
);
defparam \top/processor/sha_core/n3515_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s132  (
	.I0(\top/processor/sha_core/n3887_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_117 ),
	.I3(\top/processor/sha_core/n3515_150 ),
	.F(\top/processor/sha_core/n3887_101 )
);
defparam \top/processor/sha_core/n3887_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s181  (
	.I0(\top/processor/sha_core/n3515_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_152 ),
	.I3(\top/processor/sha_core/n3515_153 ),
	.F(\top/processor/sha_core/n3515_135 )
);
defparam \top/processor/sha_core/n3515_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s133  (
	.I0(\top/processor/sha_core/n3887_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_119 ),
	.I3(\top/processor/sha_core/n3515_153 ),
	.F(\top/processor/sha_core/n3887_103 )
);
defparam \top/processor/sha_core/n3887_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s182  (
	.I0(\top/processor/sha_core/n3515_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_155 ),
	.I3(\top/processor/sha_core/n3515_156 ),
	.F(\top/processor/sha_core/n3515_137 )
);
defparam \top/processor/sha_core/n3515_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s134  (
	.I0(\top/processor/sha_core/n3887_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_121 ),
	.I3(\top/processor/sha_core/n3515_156 ),
	.F(\top/processor/sha_core/n3887_105 )
);
defparam \top/processor/sha_core/n3887_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s183  (
	.I0(\top/processor/sha_core/n3515_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_158 ),
	.I3(\top/processor/sha_core/n3515_159 ),
	.F(\top/processor/sha_core/n3515_139 )
);
defparam \top/processor/sha_core/n3515_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s135  (
	.I0(\top/processor/sha_core/n3887_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_123 ),
	.I3(\top/processor/sha_core/n3515_159 ),
	.F(\top/processor/sha_core/n3887_107 )
);
defparam \top/processor/sha_core/n3887_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s185  (
	.I0(\top/processor/sha_core/n3490_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_164 ),
	.I3(\top/processor/sha_core/n3490_165 ),
	.F(\top/processor/sha_core/n3490_143 )
);
defparam \top/processor/sha_core/n3490_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s137  (
	.I0(\top/processor/sha_core/n3862_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_127 ),
	.I3(\top/processor/sha_core/n3490_165 ),
	.F(\top/processor/sha_core/n3862_111 )
);
defparam \top/processor/sha_core/n3862_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s184  (
	.I0(\top/processor/sha_core/n3515_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_161 ),
	.I3(\top/processor/sha_core/n3515_162 ),
	.F(\top/processor/sha_core/n3515_141 )
);
defparam \top/processor/sha_core/n3515_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s136  (
	.I0(\top/processor/sha_core/n3887_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_125 ),
	.I3(\top/processor/sha_core/n3515_162 ),
	.F(\top/processor/sha_core/n3887_109 )
);
defparam \top/processor/sha_core/n3887_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s185  (
	.I0(\top/processor/sha_core/n3515_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_164 ),
	.I3(\top/processor/sha_core/n3515_165 ),
	.F(\top/processor/sha_core/n3515_143 )
);
defparam \top/processor/sha_core/n3515_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s137  (
	.I0(\top/processor/sha_core/n3887_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_127 ),
	.I3(\top/processor/sha_core/n3515_165 ),
	.F(\top/processor/sha_core/n3887_111 )
);
defparam \top/processor/sha_core/n3887_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s186  (
	.I0(\top/processor/sha_core/n3515_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_167 ),
	.I3(\top/processor/sha_core/n3515_168 ),
	.F(\top/processor/sha_core/n3515_145 )
);
defparam \top/processor/sha_core/n3515_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s138  (
	.I0(\top/processor/sha_core/n3887_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_129 ),
	.I3(\top/processor/sha_core/n3515_168 ),
	.F(\top/processor/sha_core/n3887_113 )
);
defparam \top/processor/sha_core/n3887_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3515_s187  (
	.I0(\top/processor/sha_core/n3515_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_170 ),
	.I3(\top/processor/sha_core/n3515_171 ),
	.F(\top/processor/sha_core/n3515_147 )
);
defparam \top/processor/sha_core/n3515_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3887_s139  (
	.I0(\top/processor/sha_core/n3887_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3887_131 ),
	.I3(\top/processor/sha_core/n3515_171 ),
	.F(\top/processor/sha_core/n3887_115 )
);
defparam \top/processor/sha_core/n3887_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s180  (
	.I0(\top/processor/sha_core/n3516_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_149 ),
	.I3(\top/processor/sha_core/n3516_150 ),
	.F(\top/processor/sha_core/n3516_133 )
);
defparam \top/processor/sha_core/n3516_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s132  (
	.I0(\top/processor/sha_core/n3888_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_117 ),
	.I3(\top/processor/sha_core/n3516_150 ),
	.F(\top/processor/sha_core/n3888_101 )
);
defparam \top/processor/sha_core/n3888_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s181  (
	.I0(\top/processor/sha_core/n3516_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_152 ),
	.I3(\top/processor/sha_core/n3516_153 ),
	.F(\top/processor/sha_core/n3516_135 )
);
defparam \top/processor/sha_core/n3516_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s133  (
	.I0(\top/processor/sha_core/n3888_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_119 ),
	.I3(\top/processor/sha_core/n3516_153 ),
	.F(\top/processor/sha_core/n3888_103 )
);
defparam \top/processor/sha_core/n3888_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s182  (
	.I0(\top/processor/sha_core/n3516_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_155 ),
	.I3(\top/processor/sha_core/n3516_156 ),
	.F(\top/processor/sha_core/n3516_137 )
);
defparam \top/processor/sha_core/n3516_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s134  (
	.I0(\top/processor/sha_core/n3888_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_121 ),
	.I3(\top/processor/sha_core/n3516_156 ),
	.F(\top/processor/sha_core/n3888_105 )
);
defparam \top/processor/sha_core/n3888_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s183  (
	.I0(\top/processor/sha_core/n3516_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_158 ),
	.I3(\top/processor/sha_core/n3516_159 ),
	.F(\top/processor/sha_core/n3516_139 )
);
defparam \top/processor/sha_core/n3516_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s135  (
	.I0(\top/processor/sha_core/n3888_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_123 ),
	.I3(\top/processor/sha_core/n3516_159 ),
	.F(\top/processor/sha_core/n3888_107 )
);
defparam \top/processor/sha_core/n3888_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s184  (
	.I0(\top/processor/sha_core/n3516_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_161 ),
	.I3(\top/processor/sha_core/n3516_162 ),
	.F(\top/processor/sha_core/n3516_141 )
);
defparam \top/processor/sha_core/n3516_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s136  (
	.I0(\top/processor/sha_core/n3888_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_125 ),
	.I3(\top/processor/sha_core/n3516_162 ),
	.F(\top/processor/sha_core/n3888_109 )
);
defparam \top/processor/sha_core/n3888_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s185  (
	.I0(\top/processor/sha_core/n3516_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_164 ),
	.I3(\top/processor/sha_core/n3516_165 ),
	.F(\top/processor/sha_core/n3516_143 )
);
defparam \top/processor/sha_core/n3516_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s137  (
	.I0(\top/processor/sha_core/n3888_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_127 ),
	.I3(\top/processor/sha_core/n3516_165 ),
	.F(\top/processor/sha_core/n3888_111 )
);
defparam \top/processor/sha_core/n3888_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s186  (
	.I0(\top/processor/sha_core/n3490_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_167 ),
	.I3(\top/processor/sha_core/n3490_168 ),
	.F(\top/processor/sha_core/n3490_145 )
);
defparam \top/processor/sha_core/n3490_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s138  (
	.I0(\top/processor/sha_core/n3862_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_129 ),
	.I3(\top/processor/sha_core/n3490_168 ),
	.F(\top/processor/sha_core/n3862_113 )
);
defparam \top/processor/sha_core/n3862_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s186  (
	.I0(\top/processor/sha_core/n3516_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_167 ),
	.I3(\top/processor/sha_core/n3516_168 ),
	.F(\top/processor/sha_core/n3516_145 )
);
defparam \top/processor/sha_core/n3516_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s138  (
	.I0(\top/processor/sha_core/n3888_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_129 ),
	.I3(\top/processor/sha_core/n3516_168 ),
	.F(\top/processor/sha_core/n3888_113 )
);
defparam \top/processor/sha_core/n3888_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3516_s187  (
	.I0(\top/processor/sha_core/n3516_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_170 ),
	.I3(\top/processor/sha_core/n3516_171 ),
	.F(\top/processor/sha_core/n3516_147 )
);
defparam \top/processor/sha_core/n3516_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3888_s139  (
	.I0(\top/processor/sha_core/n3888_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3888_131 ),
	.I3(\top/processor/sha_core/n3516_171 ),
	.F(\top/processor/sha_core/n3888_115 )
);
defparam \top/processor/sha_core/n3888_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s180  (
	.I0(\top/processor/sha_core/n3517_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_149 ),
	.I3(\top/processor/sha_core/n3517_150 ),
	.F(\top/processor/sha_core/n3517_133 )
);
defparam \top/processor/sha_core/n3517_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s132  (
	.I0(\top/processor/sha_core/n3889_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_117 ),
	.I3(\top/processor/sha_core/n3517_150 ),
	.F(\top/processor/sha_core/n3889_101 )
);
defparam \top/processor/sha_core/n3889_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s181  (
	.I0(\top/processor/sha_core/n3517_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_152 ),
	.I3(\top/processor/sha_core/n3517_153 ),
	.F(\top/processor/sha_core/n3517_135 )
);
defparam \top/processor/sha_core/n3517_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s133  (
	.I0(\top/processor/sha_core/n3889_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_119 ),
	.I3(\top/processor/sha_core/n3517_153 ),
	.F(\top/processor/sha_core/n3889_103 )
);
defparam \top/processor/sha_core/n3889_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s182  (
	.I0(\top/processor/sha_core/n3517_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_155 ),
	.I3(\top/processor/sha_core/n3517_156 ),
	.F(\top/processor/sha_core/n3517_137 )
);
defparam \top/processor/sha_core/n3517_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s134  (
	.I0(\top/processor/sha_core/n3889_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_121 ),
	.I3(\top/processor/sha_core/n3517_156 ),
	.F(\top/processor/sha_core/n3889_105 )
);
defparam \top/processor/sha_core/n3889_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s183  (
	.I0(\top/processor/sha_core/n3517_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_158 ),
	.I3(\top/processor/sha_core/n3517_159 ),
	.F(\top/processor/sha_core/n3517_139 )
);
defparam \top/processor/sha_core/n3517_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s135  (
	.I0(\top/processor/sha_core/n3889_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_123 ),
	.I3(\top/processor/sha_core/n3517_159 ),
	.F(\top/processor/sha_core/n3889_107 )
);
defparam \top/processor/sha_core/n3889_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s184  (
	.I0(\top/processor/sha_core/n3517_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_161 ),
	.I3(\top/processor/sha_core/n3517_162 ),
	.F(\top/processor/sha_core/n3517_141 )
);
defparam \top/processor/sha_core/n3517_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s136  (
	.I0(\top/processor/sha_core/n3889_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_125 ),
	.I3(\top/processor/sha_core/n3517_162 ),
	.F(\top/processor/sha_core/n3889_109 )
);
defparam \top/processor/sha_core/n3889_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s185  (
	.I0(\top/processor/sha_core/n3517_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_164 ),
	.I3(\top/processor/sha_core/n3517_165 ),
	.F(\top/processor/sha_core/n3517_143 )
);
defparam \top/processor/sha_core/n3517_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s137  (
	.I0(\top/processor/sha_core/n3889_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_127 ),
	.I3(\top/processor/sha_core/n3517_165 ),
	.F(\top/processor/sha_core/n3889_111 )
);
defparam \top/processor/sha_core/n3889_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s186  (
	.I0(\top/processor/sha_core/n3517_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_167 ),
	.I3(\top/processor/sha_core/n3517_168 ),
	.F(\top/processor/sha_core/n3517_145 )
);
defparam \top/processor/sha_core/n3517_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s138  (
	.I0(\top/processor/sha_core/n3889_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_129 ),
	.I3(\top/processor/sha_core/n3517_168 ),
	.F(\top/processor/sha_core/n3889_113 )
);
defparam \top/processor/sha_core/n3889_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3517_s187  (
	.I0(\top/processor/sha_core/n3517_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_170 ),
	.I3(\top/processor/sha_core/n3517_171 ),
	.F(\top/processor/sha_core/n3517_147 )
);
defparam \top/processor/sha_core/n3517_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3889_s139  (
	.I0(\top/processor/sha_core/n3889_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3889_131 ),
	.I3(\top/processor/sha_core/n3517_171 ),
	.F(\top/processor/sha_core/n3889_115 )
);
defparam \top/processor/sha_core/n3889_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3490_s187  (
	.I0(\top/processor/sha_core/n3490_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_170 ),
	.I3(\top/processor/sha_core/n3490_171 ),
	.F(\top/processor/sha_core/n3490_147 )
);
defparam \top/processor/sha_core/n3490_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3862_s139  (
	.I0(\top/processor/sha_core/n3862_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3862_131 ),
	.I3(\top/processor/sha_core/n3490_171 ),
	.F(\top/processor/sha_core/n3862_115 )
);
defparam \top/processor/sha_core/n3862_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s180  (
	.I0(\top/processor/sha_core/n3518_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_149 ),
	.I3(\top/processor/sha_core/n3518_150 ),
	.F(\top/processor/sha_core/n3518_133 )
);
defparam \top/processor/sha_core/n3518_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s132  (
	.I0(\top/processor/sha_core/n3890_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_117 ),
	.I3(\top/processor/sha_core/n3518_150 ),
	.F(\top/processor/sha_core/n3890_101 )
);
defparam \top/processor/sha_core/n3890_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s181  (
	.I0(\top/processor/sha_core/n3518_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_152 ),
	.I3(\top/processor/sha_core/n3518_153 ),
	.F(\top/processor/sha_core/n3518_135 )
);
defparam \top/processor/sha_core/n3518_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s133  (
	.I0(\top/processor/sha_core/n3890_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_119 ),
	.I3(\top/processor/sha_core/n3518_153 ),
	.F(\top/processor/sha_core/n3890_103 )
);
defparam \top/processor/sha_core/n3890_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s182  (
	.I0(\top/processor/sha_core/n3518_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_155 ),
	.I3(\top/processor/sha_core/n3518_156 ),
	.F(\top/processor/sha_core/n3518_137 )
);
defparam \top/processor/sha_core/n3518_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s134  (
	.I0(\top/processor/sha_core/n3890_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_121 ),
	.I3(\top/processor/sha_core/n3518_156 ),
	.F(\top/processor/sha_core/n3890_105 )
);
defparam \top/processor/sha_core/n3890_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s183  (
	.I0(\top/processor/sha_core/n3518_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_158 ),
	.I3(\top/processor/sha_core/n3518_159 ),
	.F(\top/processor/sha_core/n3518_139 )
);
defparam \top/processor/sha_core/n3518_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s135  (
	.I0(\top/processor/sha_core/n3890_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_123 ),
	.I3(\top/processor/sha_core/n3518_159 ),
	.F(\top/processor/sha_core/n3890_107 )
);
defparam \top/processor/sha_core/n3890_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s184  (
	.I0(\top/processor/sha_core/n3518_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_161 ),
	.I3(\top/processor/sha_core/n3518_162 ),
	.F(\top/processor/sha_core/n3518_141 )
);
defparam \top/processor/sha_core/n3518_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s136  (
	.I0(\top/processor/sha_core/n3890_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_125 ),
	.I3(\top/processor/sha_core/n3518_162 ),
	.F(\top/processor/sha_core/n3890_109 )
);
defparam \top/processor/sha_core/n3890_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s185  (
	.I0(\top/processor/sha_core/n3518_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_164 ),
	.I3(\top/processor/sha_core/n3518_165 ),
	.F(\top/processor/sha_core/n3518_143 )
);
defparam \top/processor/sha_core/n3518_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s137  (
	.I0(\top/processor/sha_core/n3890_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_127 ),
	.I3(\top/processor/sha_core/n3518_165 ),
	.F(\top/processor/sha_core/n3890_111 )
);
defparam \top/processor/sha_core/n3890_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s186  (
	.I0(\top/processor/sha_core/n3518_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_167 ),
	.I3(\top/processor/sha_core/n3518_168 ),
	.F(\top/processor/sha_core/n3518_145 )
);
defparam \top/processor/sha_core/n3518_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s138  (
	.I0(\top/processor/sha_core/n3890_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_129 ),
	.I3(\top/processor/sha_core/n3518_168 ),
	.F(\top/processor/sha_core/n3890_113 )
);
defparam \top/processor/sha_core/n3890_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3518_s187  (
	.I0(\top/processor/sha_core/n3518_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_170 ),
	.I3(\top/processor/sha_core/n3518_171 ),
	.F(\top/processor/sha_core/n3518_147 )
);
defparam \top/processor/sha_core/n3518_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3890_s139  (
	.I0(\top/processor/sha_core/n3890_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3890_131 ),
	.I3(\top/processor/sha_core/n3518_171 ),
	.F(\top/processor/sha_core/n3890_115 )
);
defparam \top/processor/sha_core/n3890_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s180  (
	.I0(\top/processor/sha_core/n3519_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_149 ),
	.I3(\top/processor/sha_core/n3519_150 ),
	.F(\top/processor/sha_core/n3519_133 )
);
defparam \top/processor/sha_core/n3519_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s132  (
	.I0(\top/processor/sha_core/n3891_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_117 ),
	.I3(\top/processor/sha_core/n3519_150 ),
	.F(\top/processor/sha_core/n3891_101 )
);
defparam \top/processor/sha_core/n3891_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s181  (
	.I0(\top/processor/sha_core/n3519_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_152 ),
	.I3(\top/processor/sha_core/n3519_153 ),
	.F(\top/processor/sha_core/n3519_135 )
);
defparam \top/processor/sha_core/n3519_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s133  (
	.I0(\top/processor/sha_core/n3891_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_119 ),
	.I3(\top/processor/sha_core/n3519_153 ),
	.F(\top/processor/sha_core/n3891_103 )
);
defparam \top/processor/sha_core/n3891_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3491_s180  (
	.I0(\top/processor/sha_core/n3491_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_149 ),
	.I3(\top/processor/sha_core/n3491_150 ),
	.F(\top/processor/sha_core/n3491_133 )
);
defparam \top/processor/sha_core/n3491_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s132  (
	.I0(\top/processor/sha_core/n3863_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_117 ),
	.I3(\top/processor/sha_core/n3491_150 ),
	.F(\top/processor/sha_core/n3863_101 )
);
defparam \top/processor/sha_core/n3863_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s182  (
	.I0(\top/processor/sha_core/n3519_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_155 ),
	.I3(\top/processor/sha_core/n3519_156 ),
	.F(\top/processor/sha_core/n3519_137 )
);
defparam \top/processor/sha_core/n3519_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s134  (
	.I0(\top/processor/sha_core/n3891_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_121 ),
	.I3(\top/processor/sha_core/n3519_156 ),
	.F(\top/processor/sha_core/n3891_105 )
);
defparam \top/processor/sha_core/n3891_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s183  (
	.I0(\top/processor/sha_core/n3519_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_158 ),
	.I3(\top/processor/sha_core/n3519_159 ),
	.F(\top/processor/sha_core/n3519_139 )
);
defparam \top/processor/sha_core/n3519_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s135  (
	.I0(\top/processor/sha_core/n3891_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_123 ),
	.I3(\top/processor/sha_core/n3519_159 ),
	.F(\top/processor/sha_core/n3891_107 )
);
defparam \top/processor/sha_core/n3891_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s184  (
	.I0(\top/processor/sha_core/n3519_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_161 ),
	.I3(\top/processor/sha_core/n3519_162 ),
	.F(\top/processor/sha_core/n3519_141 )
);
defparam \top/processor/sha_core/n3519_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s136  (
	.I0(\top/processor/sha_core/n3891_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_125 ),
	.I3(\top/processor/sha_core/n3519_162 ),
	.F(\top/processor/sha_core/n3891_109 )
);
defparam \top/processor/sha_core/n3891_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s185  (
	.I0(\top/processor/sha_core/n3519_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_164 ),
	.I3(\top/processor/sha_core/n3519_165 ),
	.F(\top/processor/sha_core/n3519_143 )
);
defparam \top/processor/sha_core/n3519_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s137  (
	.I0(\top/processor/sha_core/n3891_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_127 ),
	.I3(\top/processor/sha_core/n3519_165 ),
	.F(\top/processor/sha_core/n3891_111 )
);
defparam \top/processor/sha_core/n3891_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s186  (
	.I0(\top/processor/sha_core/n3519_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_167 ),
	.I3(\top/processor/sha_core/n3519_168 ),
	.F(\top/processor/sha_core/n3519_145 )
);
defparam \top/processor/sha_core/n3519_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s138  (
	.I0(\top/processor/sha_core/n3891_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_129 ),
	.I3(\top/processor/sha_core/n3519_168 ),
	.F(\top/processor/sha_core/n3891_113 )
);
defparam \top/processor/sha_core/n3891_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3519_s187  (
	.I0(\top/processor/sha_core/n3519_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_170 ),
	.I3(\top/processor/sha_core/n3519_171 ),
	.F(\top/processor/sha_core/n3519_147 )
);
defparam \top/processor/sha_core/n3519_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3891_s139  (
	.I0(\top/processor/sha_core/n3891_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3891_131 ),
	.I3(\top/processor/sha_core/n3519_171 ),
	.F(\top/processor/sha_core/n3891_115 )
);
defparam \top/processor/sha_core/n3891_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s135  (
	.I0(\top/processor/sha_core/n3607_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [31]),
	.I3(\top/processor/sha_core/w[0] [31]),
	.F(\top/processor/sha_core/n3607_149 )
);
defparam \top/processor/sha_core/n3705_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s135  (
	.I0(\top/processor/sha_core/n3608_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [30]),
	.I3(\top/processor/sha_core/w[0] [30]),
	.F(\top/processor/sha_core/n3608_149 )
);
defparam \top/processor/sha_core/n3706_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s135  (
	.I0(\top/processor/sha_core/n3609_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [29]),
	.I3(\top/processor/sha_core/w[0] [29]),
	.F(\top/processor/sha_core/n3609_149 )
);
defparam \top/processor/sha_core/n3707_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s135  (
	.I0(\top/processor/sha_core/n3610_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [28]),
	.I3(\top/processor/sha_core/w[0] [28]),
	.F(\top/processor/sha_core/n3610_149 )
);
defparam \top/processor/sha_core/n3708_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s135  (
	.I0(\top/processor/sha_core/n3611_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [27]),
	.I3(\top/processor/sha_core/w[0] [27]),
	.F(\top/processor/sha_core/n3611_149 )
);
defparam \top/processor/sha_core/n3709_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s135  (
	.I0(\top/processor/sha_core/n3612_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [26]),
	.I3(\top/processor/sha_core/w[0] [26]),
	.F(\top/processor/sha_core/n3612_149 )
);
defparam \top/processor/sha_core/n3710_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s135  (
	.I0(\top/processor/sha_core/n3613_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [25]),
	.I3(\top/processor/sha_core/w[0] [25]),
	.F(\top/processor/sha_core/n3613_149 )
);
defparam \top/processor/sha_core/n3711_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3491_s181  (
	.I0(\top/processor/sha_core/n3491_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_152 ),
	.I3(\top/processor/sha_core/n3491_153 ),
	.F(\top/processor/sha_core/n3491_135 )
);
defparam \top/processor/sha_core/n3491_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s133  (
	.I0(\top/processor/sha_core/n3863_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_119 ),
	.I3(\top/processor/sha_core/n3491_153 ),
	.F(\top/processor/sha_core/n3863_103 )
);
defparam \top/processor/sha_core/n3863_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3712_s135  (
	.I0(\top/processor/sha_core/n3614_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [24]),
	.I3(\top/processor/sha_core/w[0] [24]),
	.F(\top/processor/sha_core/n3614_149 )
);
defparam \top/processor/sha_core/n3712_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s135  (
	.I0(\top/processor/sha_core/n3615_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [23]),
	.I3(\top/processor/sha_core/w[0] [23]),
	.F(\top/processor/sha_core/n3615_149 )
);
defparam \top/processor/sha_core/n3713_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s135  (
	.I0(\top/processor/sha_core/n3616_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [22]),
	.I3(\top/processor/sha_core/w[0] [22]),
	.F(\top/processor/sha_core/n3616_149 )
);
defparam \top/processor/sha_core/n3714_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s135  (
	.I0(\top/processor/sha_core/n3617_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [21]),
	.I3(\top/processor/sha_core/w[0] [21]),
	.F(\top/processor/sha_core/n3617_149 )
);
defparam \top/processor/sha_core/n3715_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s135  (
	.I0(\top/processor/sha_core/n3618_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [20]),
	.I3(\top/processor/sha_core/w[0] [20]),
	.F(\top/processor/sha_core/n3618_149 )
);
defparam \top/processor/sha_core/n3716_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s135  (
	.I0(\top/processor/sha_core/n3619_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [19]),
	.I3(\top/processor/sha_core/w[0] [19]),
	.F(\top/processor/sha_core/n3619_149 )
);
defparam \top/processor/sha_core/n3717_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s135  (
	.I0(\top/processor/sha_core/n3620_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [18]),
	.I3(\top/processor/sha_core/w[0] [18]),
	.F(\top/processor/sha_core/n3620_149 )
);
defparam \top/processor/sha_core/n3718_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s135  (
	.I0(\top/processor/sha_core/n3621_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [17]),
	.I3(\top/processor/sha_core/w[0] [17]),
	.F(\top/processor/sha_core/n3621_149 )
);
defparam \top/processor/sha_core/n3719_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s135  (
	.I0(\top/processor/sha_core/n3622_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [16]),
	.I3(\top/processor/sha_core/w[0] [16]),
	.F(\top/processor/sha_core/n3622_149 )
);
defparam \top/processor/sha_core/n3720_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s135  (
	.I0(\top/processor/sha_core/n3623_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [15]),
	.I3(\top/processor/sha_core/w[0] [15]),
	.F(\top/processor/sha_core/n3623_149 )
);
defparam \top/processor/sha_core/n3721_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s135  (
	.I0(\top/processor/sha_core/n3624_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [14]),
	.I3(\top/processor/sha_core/w[0] [14]),
	.F(\top/processor/sha_core/n3624_149 )
);
defparam \top/processor/sha_core/n3722_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s135  (
	.I0(\top/processor/sha_core/n3625_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [13]),
	.I3(\top/processor/sha_core/w[0] [13]),
	.F(\top/processor/sha_core/n3625_149 )
);
defparam \top/processor/sha_core/n3723_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s135  (
	.I0(\top/processor/sha_core/n3626_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [12]),
	.I3(\top/processor/sha_core/w[0] [12]),
	.F(\top/processor/sha_core/n3626_149 )
);
defparam \top/processor/sha_core/n3724_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s135  (
	.I0(\top/processor/sha_core/n3627_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [11]),
	.I3(\top/processor/sha_core/w[0] [11]),
	.F(\top/processor/sha_core/n3627_149 )
);
defparam \top/processor/sha_core/n3725_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s135  (
	.I0(\top/processor/sha_core/n3628_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [10]),
	.I3(\top/processor/sha_core/w[0] [10]),
	.F(\top/processor/sha_core/n3628_149 )
);
defparam \top/processor/sha_core/n3726_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s135  (
	.I0(\top/processor/sha_core/n3629_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [9]),
	.I3(\top/processor/sha_core/w[0] [9]),
	.F(\top/processor/sha_core/n3629_149 )
);
defparam \top/processor/sha_core/n3727_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s135  (
	.I0(\top/processor/sha_core/n3630_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [8]),
	.I3(\top/processor/sha_core/w[0] [8]),
	.F(\top/processor/sha_core/n3630_149 )
);
defparam \top/processor/sha_core/n3728_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s135  (
	.I0(\top/processor/sha_core/n3631_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [7]),
	.I3(\top/processor/sha_core/w[0] [7]),
	.F(\top/processor/sha_core/n3631_149 )
);
defparam \top/processor/sha_core/n3729_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s135  (
	.I0(\top/processor/sha_core/n3632_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [6]),
	.I3(\top/processor/sha_core/w[0] [6]),
	.F(\top/processor/sha_core/n3632_149 )
);
defparam \top/processor/sha_core/n3730_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s135  (
	.I0(\top/processor/sha_core/n3633_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [5]),
	.I3(\top/processor/sha_core/w[0] [5]),
	.F(\top/processor/sha_core/n3633_149 )
);
defparam \top/processor/sha_core/n3731_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3491_s182  (
	.I0(\top/processor/sha_core/n3491_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_155 ),
	.I3(\top/processor/sha_core/n3491_156 ),
	.F(\top/processor/sha_core/n3491_137 )
);
defparam \top/processor/sha_core/n3491_s182 .INIT=16'hD951;
LUT4 \top/processor/sha_core/n3863_s134  (
	.I0(\top/processor/sha_core/n3863_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_121 ),
	.I3(\top/processor/sha_core/n3491_156 ),
	.F(\top/processor/sha_core/n3863_105 )
);
defparam \top/processor/sha_core/n3863_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3732_s135  (
	.I0(\top/processor/sha_core/n3634_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [4]),
	.I3(\top/processor/sha_core/w[0] [4]),
	.F(\top/processor/sha_core/n3634_149 )
);
defparam \top/processor/sha_core/n3732_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s135  (
	.I0(\top/processor/sha_core/n3635_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [3]),
	.I3(\top/processor/sha_core/w[0] [3]),
	.F(\top/processor/sha_core/n3635_149 )
);
defparam \top/processor/sha_core/n3733_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s135  (
	.I0(\top/processor/sha_core/n3636_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [2]),
	.I3(\top/processor/sha_core/w[0] [2]),
	.F(\top/processor/sha_core/n3636_149 )
);
defparam \top/processor/sha_core/n3734_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s135  (
	.I0(\top/processor/sha_core/n3637_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [1]),
	.I3(\top/processor/sha_core/w[0] [1]),
	.F(\top/processor/sha_core/n3637_149 )
);
defparam \top/processor/sha_core/n3735_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s135  (
	.I0(\top/processor/sha_core/n3638_172 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[2] [0]),
	.I3(\top/processor/sha_core/w[0] [0]),
	.F(\top/processor/sha_core/n3638_149 )
);
defparam \top/processor/sha_core/n3736_s135 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3491_s183  (
	.I0(\top/processor/sha_core/n3491_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_158 ),
	.I3(\top/processor/sha_core/n3491_159 ),
	.F(\top/processor/sha_core/n3491_139 )
);
defparam \top/processor/sha_core/n3491_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s135  (
	.I0(\top/processor/sha_core/n3863_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_123 ),
	.I3(\top/processor/sha_core/n3491_159 ),
	.F(\top/processor/sha_core/n3863_107 )
);
defparam \top/processor/sha_core/n3863_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s136  (
	.I0(\top/processor/sha_core/n3607_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [31]),
	.I3(\top/processor/sha_core/w[4] [31]),
	.F(\top/processor/sha_core/n3607_151 )
);
defparam \top/processor/sha_core/n3705_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s136  (
	.I0(\top/processor/sha_core/n3608_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [30]),
	.I3(\top/processor/sha_core/w[4] [30]),
	.F(\top/processor/sha_core/n3608_151 )
);
defparam \top/processor/sha_core/n3706_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s136  (
	.I0(\top/processor/sha_core/n3609_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [29]),
	.I3(\top/processor/sha_core/w[4] [29]),
	.F(\top/processor/sha_core/n3609_151 )
);
defparam \top/processor/sha_core/n3707_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3491_s184  (
	.I0(\top/processor/sha_core/n3491_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_161 ),
	.I3(\top/processor/sha_core/n3491_162 ),
	.F(\top/processor/sha_core/n3491_141 )
);
defparam \top/processor/sha_core/n3491_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s136  (
	.I0(\top/processor/sha_core/n3863_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_125 ),
	.I3(\top/processor/sha_core/n3491_162 ),
	.F(\top/processor/sha_core/n3863_109 )
);
defparam \top/processor/sha_core/n3863_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3708_s136  (
	.I0(\top/processor/sha_core/n3610_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [28]),
	.I3(\top/processor/sha_core/w[4] [28]),
	.F(\top/processor/sha_core/n3610_151 )
);
defparam \top/processor/sha_core/n3708_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s136  (
	.I0(\top/processor/sha_core/n3611_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [27]),
	.I3(\top/processor/sha_core/w[4] [27]),
	.F(\top/processor/sha_core/n3611_151 )
);
defparam \top/processor/sha_core/n3709_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s136  (
	.I0(\top/processor/sha_core/n3612_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [26]),
	.I3(\top/processor/sha_core/w[4] [26]),
	.F(\top/processor/sha_core/n3612_151 )
);
defparam \top/processor/sha_core/n3710_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s136  (
	.I0(\top/processor/sha_core/n3613_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [25]),
	.I3(\top/processor/sha_core/w[4] [25]),
	.F(\top/processor/sha_core/n3613_151 )
);
defparam \top/processor/sha_core/n3711_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s136  (
	.I0(\top/processor/sha_core/n3614_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [24]),
	.I3(\top/processor/sha_core/w[4] [24]),
	.F(\top/processor/sha_core/n3614_151 )
);
defparam \top/processor/sha_core/n3712_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s136  (
	.I0(\top/processor/sha_core/n3615_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [23]),
	.I3(\top/processor/sha_core/w[4] [23]),
	.F(\top/processor/sha_core/n3615_151 )
);
defparam \top/processor/sha_core/n3713_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s136  (
	.I0(\top/processor/sha_core/n3616_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [22]),
	.I3(\top/processor/sha_core/w[4] [22]),
	.F(\top/processor/sha_core/n3616_151 )
);
defparam \top/processor/sha_core/n3714_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s136  (
	.I0(\top/processor/sha_core/n3617_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [21]),
	.I3(\top/processor/sha_core/w[4] [21]),
	.F(\top/processor/sha_core/n3617_151 )
);
defparam \top/processor/sha_core/n3715_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s136  (
	.I0(\top/processor/sha_core/n3618_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [20]),
	.I3(\top/processor/sha_core/w[4] [20]),
	.F(\top/processor/sha_core/n3618_151 )
);
defparam \top/processor/sha_core/n3716_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s136  (
	.I0(\top/processor/sha_core/n3619_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [19]),
	.I3(\top/processor/sha_core/w[4] [19]),
	.F(\top/processor/sha_core/n3619_151 )
);
defparam \top/processor/sha_core/n3717_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s136  (
	.I0(\top/processor/sha_core/n3620_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [18]),
	.I3(\top/processor/sha_core/w[4] [18]),
	.F(\top/processor/sha_core/n3620_151 )
);
defparam \top/processor/sha_core/n3718_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s136  (
	.I0(\top/processor/sha_core/n3621_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [17]),
	.I3(\top/processor/sha_core/w[4] [17]),
	.F(\top/processor/sha_core/n3621_151 )
);
defparam \top/processor/sha_core/n3719_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s136  (
	.I0(\top/processor/sha_core/n3622_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [16]),
	.I3(\top/processor/sha_core/w[4] [16]),
	.F(\top/processor/sha_core/n3622_151 )
);
defparam \top/processor/sha_core/n3720_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s136  (
	.I0(\top/processor/sha_core/n3623_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [15]),
	.I3(\top/processor/sha_core/w[4] [15]),
	.F(\top/processor/sha_core/n3623_151 )
);
defparam \top/processor/sha_core/n3721_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s136  (
	.I0(\top/processor/sha_core/n3624_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [14]),
	.I3(\top/processor/sha_core/w[4] [14]),
	.F(\top/processor/sha_core/n3624_151 )
);
defparam \top/processor/sha_core/n3722_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s136  (
	.I0(\top/processor/sha_core/n3625_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [13]),
	.I3(\top/processor/sha_core/w[4] [13]),
	.F(\top/processor/sha_core/n3625_151 )
);
defparam \top/processor/sha_core/n3723_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s136  (
	.I0(\top/processor/sha_core/n3626_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [12]),
	.I3(\top/processor/sha_core/w[4] [12]),
	.F(\top/processor/sha_core/n3626_151 )
);
defparam \top/processor/sha_core/n3724_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s136  (
	.I0(\top/processor/sha_core/n3627_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [11]),
	.I3(\top/processor/sha_core/w[4] [11]),
	.F(\top/processor/sha_core/n3627_151 )
);
defparam \top/processor/sha_core/n3725_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s136  (
	.I0(\top/processor/sha_core/n3628_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [10]),
	.I3(\top/processor/sha_core/w[4] [10]),
	.F(\top/processor/sha_core/n3628_151 )
);
defparam \top/processor/sha_core/n3726_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s136  (
	.I0(\top/processor/sha_core/n3629_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [9]),
	.I3(\top/processor/sha_core/w[4] [9]),
	.F(\top/processor/sha_core/n3629_151 )
);
defparam \top/processor/sha_core/n3727_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3491_s185  (
	.I0(\top/processor/sha_core/n3491_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_164 ),
	.I3(\top/processor/sha_core/n3491_165 ),
	.F(\top/processor/sha_core/n3491_143 )
);
defparam \top/processor/sha_core/n3491_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s137  (
	.I0(\top/processor/sha_core/n3863_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_127 ),
	.I3(\top/processor/sha_core/n3491_165 ),
	.F(\top/processor/sha_core/n3863_111 )
);
defparam \top/processor/sha_core/n3863_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s182  (
	.I0(\top/processor/sha_core/n3488_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_164 ),
	.I3(\top/processor/sha_core/n3488_165 ),
	.F(\top/processor/sha_core/n3488_143 )
);
defparam \top/processor/sha_core/n3488_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s134  (
	.I0(\top/processor/sha_core/n3860_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_127 ),
	.I3(\top/processor/sha_core/n3488_165 ),
	.F(\top/processor/sha_core/n3860_111 )
);
defparam \top/processor/sha_core/n3860_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3728_s136  (
	.I0(\top/processor/sha_core/n3630_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [8]),
	.I3(\top/processor/sha_core/w[4] [8]),
	.F(\top/processor/sha_core/n3630_151 )
);
defparam \top/processor/sha_core/n3728_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s136  (
	.I0(\top/processor/sha_core/n3631_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [7]),
	.I3(\top/processor/sha_core/w[4] [7]),
	.F(\top/processor/sha_core/n3631_151 )
);
defparam \top/processor/sha_core/n3729_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s136  (
	.I0(\top/processor/sha_core/n3632_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [6]),
	.I3(\top/processor/sha_core/w[4] [6]),
	.F(\top/processor/sha_core/n3632_151 )
);
defparam \top/processor/sha_core/n3730_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s136  (
	.I0(\top/processor/sha_core/n3633_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [5]),
	.I3(\top/processor/sha_core/w[4] [5]),
	.F(\top/processor/sha_core/n3633_151 )
);
defparam \top/processor/sha_core/n3731_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s136  (
	.I0(\top/processor/sha_core/n3634_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [4]),
	.I3(\top/processor/sha_core/w[4] [4]),
	.F(\top/processor/sha_core/n3634_151 )
);
defparam \top/processor/sha_core/n3732_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s136  (
	.I0(\top/processor/sha_core/n3635_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [3]),
	.I3(\top/processor/sha_core/w[4] [3]),
	.F(\top/processor/sha_core/n3635_151 )
);
defparam \top/processor/sha_core/n3733_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s136  (
	.I0(\top/processor/sha_core/n3636_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [2]),
	.I3(\top/processor/sha_core/w[4] [2]),
	.F(\top/processor/sha_core/n3636_151 )
);
defparam \top/processor/sha_core/n3734_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s136  (
	.I0(\top/processor/sha_core/n3637_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [1]),
	.I3(\top/processor/sha_core/w[4] [1]),
	.F(\top/processor/sha_core/n3637_151 )
);
defparam \top/processor/sha_core/n3735_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s136  (
	.I0(\top/processor/sha_core/n3638_173 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[6] [0]),
	.I3(\top/processor/sha_core/w[4] [0]),
	.F(\top/processor/sha_core/n3638_151 )
);
defparam \top/processor/sha_core/n3736_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3491_s186  (
	.I0(\top/processor/sha_core/n3491_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_167 ),
	.I3(\top/processor/sha_core/n3491_168 ),
	.F(\top/processor/sha_core/n3491_145 )
);
defparam \top/processor/sha_core/n3491_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s138  (
	.I0(\top/processor/sha_core/n3863_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_129 ),
	.I3(\top/processor/sha_core/n3491_168 ),
	.F(\top/processor/sha_core/n3863_113 )
);
defparam \top/processor/sha_core/n3863_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3491_s187  (
	.I0(\top/processor/sha_core/n3491_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_170 ),
	.I3(\top/processor/sha_core/n3491_171 ),
	.F(\top/processor/sha_core/n3491_147 )
);
defparam \top/processor/sha_core/n3491_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3863_s139  (
	.I0(\top/processor/sha_core/n3863_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3863_131 ),
	.I3(\top/processor/sha_core/n3491_171 ),
	.F(\top/processor/sha_core/n3863_115 )
);
defparam \top/processor/sha_core/n3863_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s137  (
	.I0(\top/processor/sha_core/n3607_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [31]),
	.I3(\top/processor/sha_core/w[8] [31]),
	.F(\top/processor/sha_core/n3607_153 )
);
defparam \top/processor/sha_core/n3705_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s137  (
	.I0(\top/processor/sha_core/n3608_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [30]),
	.I3(\top/processor/sha_core/w[8] [30]),
	.F(\top/processor/sha_core/n3608_153 )
);
defparam \top/processor/sha_core/n3706_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s137  (
	.I0(\top/processor/sha_core/n3609_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [29]),
	.I3(\top/processor/sha_core/w[8] [29]),
	.F(\top/processor/sha_core/n3609_153 )
);
defparam \top/processor/sha_core/n3707_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s137  (
	.I0(\top/processor/sha_core/n3610_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [28]),
	.I3(\top/processor/sha_core/w[8] [28]),
	.F(\top/processor/sha_core/n3610_153 )
);
defparam \top/processor/sha_core/n3708_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s137  (
	.I0(\top/processor/sha_core/n3611_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [27]),
	.I3(\top/processor/sha_core/w[8] [27]),
	.F(\top/processor/sha_core/n3611_153 )
);
defparam \top/processor/sha_core/n3709_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s137  (
	.I0(\top/processor/sha_core/n3612_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [26]),
	.I3(\top/processor/sha_core/w[8] [26]),
	.F(\top/processor/sha_core/n3612_153 )
);
defparam \top/processor/sha_core/n3710_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s137  (
	.I0(\top/processor/sha_core/n3613_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [25]),
	.I3(\top/processor/sha_core/w[8] [25]),
	.F(\top/processor/sha_core/n3613_153 )
);
defparam \top/processor/sha_core/n3711_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s137  (
	.I0(\top/processor/sha_core/n3614_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [24]),
	.I3(\top/processor/sha_core/w[8] [24]),
	.F(\top/processor/sha_core/n3614_153 )
);
defparam \top/processor/sha_core/n3712_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s137  (
	.I0(\top/processor/sha_core/n3615_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [23]),
	.I3(\top/processor/sha_core/w[8] [23]),
	.F(\top/processor/sha_core/n3615_153 )
);
defparam \top/processor/sha_core/n3713_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s137  (
	.I0(\top/processor/sha_core/n3616_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [22]),
	.I3(\top/processor/sha_core/w[8] [22]),
	.F(\top/processor/sha_core/n3616_153 )
);
defparam \top/processor/sha_core/n3714_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s137  (
	.I0(\top/processor/sha_core/n3617_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [21]),
	.I3(\top/processor/sha_core/w[8] [21]),
	.F(\top/processor/sha_core/n3617_153 )
);
defparam \top/processor/sha_core/n3715_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s137  (
	.I0(\top/processor/sha_core/n3618_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [20]),
	.I3(\top/processor/sha_core/w[8] [20]),
	.F(\top/processor/sha_core/n3618_153 )
);
defparam \top/processor/sha_core/n3716_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s137  (
	.I0(\top/processor/sha_core/n3619_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [19]),
	.I3(\top/processor/sha_core/w[8] [19]),
	.F(\top/processor/sha_core/n3619_153 )
);
defparam \top/processor/sha_core/n3717_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s137  (
	.I0(\top/processor/sha_core/n3620_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [18]),
	.I3(\top/processor/sha_core/w[8] [18]),
	.F(\top/processor/sha_core/n3620_153 )
);
defparam \top/processor/sha_core/n3718_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s137  (
	.I0(\top/processor/sha_core/n3621_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [17]),
	.I3(\top/processor/sha_core/w[8] [17]),
	.F(\top/processor/sha_core/n3621_153 )
);
defparam \top/processor/sha_core/n3719_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s137  (
	.I0(\top/processor/sha_core/n3622_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [16]),
	.I3(\top/processor/sha_core/w[8] [16]),
	.F(\top/processor/sha_core/n3622_153 )
);
defparam \top/processor/sha_core/n3720_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s137  (
	.I0(\top/processor/sha_core/n3623_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [15]),
	.I3(\top/processor/sha_core/w[8] [15]),
	.F(\top/processor/sha_core/n3623_153 )
);
defparam \top/processor/sha_core/n3721_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s137  (
	.I0(\top/processor/sha_core/n3624_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [14]),
	.I3(\top/processor/sha_core/w[8] [14]),
	.F(\top/processor/sha_core/n3624_153 )
);
defparam \top/processor/sha_core/n3722_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s137  (
	.I0(\top/processor/sha_core/n3625_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [13]),
	.I3(\top/processor/sha_core/w[8] [13]),
	.F(\top/processor/sha_core/n3625_153 )
);
defparam \top/processor/sha_core/n3723_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3492_s180  (
	.I0(\top/processor/sha_core/n3492_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_149 ),
	.I3(\top/processor/sha_core/n3492_150 ),
	.F(\top/processor/sha_core/n3492_133 )
);
defparam \top/processor/sha_core/n3492_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s132  (
	.I0(\top/processor/sha_core/n3864_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_117 ),
	.I3(\top/processor/sha_core/n3492_150 ),
	.F(\top/processor/sha_core/n3864_101 )
);
defparam \top/processor/sha_core/n3864_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3724_s137  (
	.I0(\top/processor/sha_core/n3626_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [12]),
	.I3(\top/processor/sha_core/w[8] [12]),
	.F(\top/processor/sha_core/n3626_153 )
);
defparam \top/processor/sha_core/n3724_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s137  (
	.I0(\top/processor/sha_core/n3627_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [11]),
	.I3(\top/processor/sha_core/w[8] [11]),
	.F(\top/processor/sha_core/n3627_153 )
);
defparam \top/processor/sha_core/n3725_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s137  (
	.I0(\top/processor/sha_core/n3628_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [10]),
	.I3(\top/processor/sha_core/w[8] [10]),
	.F(\top/processor/sha_core/n3628_153 )
);
defparam \top/processor/sha_core/n3726_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s137  (
	.I0(\top/processor/sha_core/n3629_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [9]),
	.I3(\top/processor/sha_core/w[8] [9]),
	.F(\top/processor/sha_core/n3629_153 )
);
defparam \top/processor/sha_core/n3727_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s137  (
	.I0(\top/processor/sha_core/n3630_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [8]),
	.I3(\top/processor/sha_core/w[8] [8]),
	.F(\top/processor/sha_core/n3630_153 )
);
defparam \top/processor/sha_core/n3728_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s137  (
	.I0(\top/processor/sha_core/n3631_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [7]),
	.I3(\top/processor/sha_core/w[8] [7]),
	.F(\top/processor/sha_core/n3631_153 )
);
defparam \top/processor/sha_core/n3729_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s137  (
	.I0(\top/processor/sha_core/n3632_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [6]),
	.I3(\top/processor/sha_core/w[8] [6]),
	.F(\top/processor/sha_core/n3632_153 )
);
defparam \top/processor/sha_core/n3730_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s137  (
	.I0(\top/processor/sha_core/n3633_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [5]),
	.I3(\top/processor/sha_core/w[8] [5]),
	.F(\top/processor/sha_core/n3633_153 )
);
defparam \top/processor/sha_core/n3731_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s137  (
	.I0(\top/processor/sha_core/n3634_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [4]),
	.I3(\top/processor/sha_core/w[8] [4]),
	.F(\top/processor/sha_core/n3634_153 )
);
defparam \top/processor/sha_core/n3732_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s137  (
	.I0(\top/processor/sha_core/n3635_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [3]),
	.I3(\top/processor/sha_core/w[8] [3]),
	.F(\top/processor/sha_core/n3635_153 )
);
defparam \top/processor/sha_core/n3733_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s137  (
	.I0(\top/processor/sha_core/n3636_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [2]),
	.I3(\top/processor/sha_core/w[8] [2]),
	.F(\top/processor/sha_core/n3636_153 )
);
defparam \top/processor/sha_core/n3734_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s137  (
	.I0(\top/processor/sha_core/n3637_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [1]),
	.I3(\top/processor/sha_core/w[8] [1]),
	.F(\top/processor/sha_core/n3637_153 )
);
defparam \top/processor/sha_core/n3735_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s137  (
	.I0(\top/processor/sha_core/n3638_174 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[10] [0]),
	.I3(\top/processor/sha_core/w[8] [0]),
	.F(\top/processor/sha_core/n3638_153 )
);
defparam \top/processor/sha_core/n3736_s137 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3492_s181  (
	.I0(\top/processor/sha_core/n3492_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_152 ),
	.I3(\top/processor/sha_core/n3492_153 ),
	.F(\top/processor/sha_core/n3492_135 )
);
defparam \top/processor/sha_core/n3492_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s133  (
	.I0(\top/processor/sha_core/n3864_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_119 ),
	.I3(\top/processor/sha_core/n3492_153 ),
	.F(\top/processor/sha_core/n3864_103 )
);
defparam \top/processor/sha_core/n3864_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3492_s182  (
	.I0(\top/processor/sha_core/n3492_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_155 ),
	.I3(\top/processor/sha_core/n3492_156 ),
	.F(\top/processor/sha_core/n3492_137 )
);
defparam \top/processor/sha_core/n3492_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s134  (
	.I0(\top/processor/sha_core/n3864_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_121 ),
	.I3(\top/processor/sha_core/n3492_156 ),
	.F(\top/processor/sha_core/n3864_105 )
);
defparam \top/processor/sha_core/n3864_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s138  (
	.I0(\top/processor/sha_core/n3607_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [31]),
	.I3(\top/processor/sha_core/w[12] [31]),
	.F(\top/processor/sha_core/n3607_155 )
);
defparam \top/processor/sha_core/n3705_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s138  (
	.I0(\top/processor/sha_core/n3608_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [30]),
	.I3(\top/processor/sha_core/w[12] [30]),
	.F(\top/processor/sha_core/n3608_155 )
);
defparam \top/processor/sha_core/n3706_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s138  (
	.I0(\top/processor/sha_core/n3609_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [29]),
	.I3(\top/processor/sha_core/w[12] [29]),
	.F(\top/processor/sha_core/n3609_155 )
);
defparam \top/processor/sha_core/n3707_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s138  (
	.I0(\top/processor/sha_core/n3610_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [28]),
	.I3(\top/processor/sha_core/w[12] [28]),
	.F(\top/processor/sha_core/n3610_155 )
);
defparam \top/processor/sha_core/n3708_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s138  (
	.I0(\top/processor/sha_core/n3611_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [27]),
	.I3(\top/processor/sha_core/w[12] [27]),
	.F(\top/processor/sha_core/n3611_155 )
);
defparam \top/processor/sha_core/n3709_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s138  (
	.I0(\top/processor/sha_core/n3612_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [26]),
	.I3(\top/processor/sha_core/w[12] [26]),
	.F(\top/processor/sha_core/n3612_155 )
);
defparam \top/processor/sha_core/n3710_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s138  (
	.I0(\top/processor/sha_core/n3613_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [25]),
	.I3(\top/processor/sha_core/w[12] [25]),
	.F(\top/processor/sha_core/n3613_155 )
);
defparam \top/processor/sha_core/n3711_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s138  (
	.I0(\top/processor/sha_core/n3614_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [24]),
	.I3(\top/processor/sha_core/w[12] [24]),
	.F(\top/processor/sha_core/n3614_155 )
);
defparam \top/processor/sha_core/n3712_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s138  (
	.I0(\top/processor/sha_core/n3615_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [23]),
	.I3(\top/processor/sha_core/w[12] [23]),
	.F(\top/processor/sha_core/n3615_155 )
);
defparam \top/processor/sha_core/n3713_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s138  (
	.I0(\top/processor/sha_core/n3616_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [22]),
	.I3(\top/processor/sha_core/w[12] [22]),
	.F(\top/processor/sha_core/n3616_155 )
);
defparam \top/processor/sha_core/n3714_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s138  (
	.I0(\top/processor/sha_core/n3617_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [21]),
	.I3(\top/processor/sha_core/w[12] [21]),
	.F(\top/processor/sha_core/n3617_155 )
);
defparam \top/processor/sha_core/n3715_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s138  (
	.I0(\top/processor/sha_core/n3618_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [20]),
	.I3(\top/processor/sha_core/w[12] [20]),
	.F(\top/processor/sha_core/n3618_155 )
);
defparam \top/processor/sha_core/n3716_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s138  (
	.I0(\top/processor/sha_core/n3619_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [19]),
	.I3(\top/processor/sha_core/w[12] [19]),
	.F(\top/processor/sha_core/n3619_155 )
);
defparam \top/processor/sha_core/n3717_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s138  (
	.I0(\top/processor/sha_core/n3620_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [18]),
	.I3(\top/processor/sha_core/w[12] [18]),
	.F(\top/processor/sha_core/n3620_155 )
);
defparam \top/processor/sha_core/n3718_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s138  (
	.I0(\top/processor/sha_core/n3621_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [17]),
	.I3(\top/processor/sha_core/w[12] [17]),
	.F(\top/processor/sha_core/n3621_155 )
);
defparam \top/processor/sha_core/n3719_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3492_s183  (
	.I0(\top/processor/sha_core/n3492_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_158 ),
	.I3(\top/processor/sha_core/n3492_159 ),
	.F(\top/processor/sha_core/n3492_139 )
);
defparam \top/processor/sha_core/n3492_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s135  (
	.I0(\top/processor/sha_core/n3864_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_123 ),
	.I3(\top/processor/sha_core/n3492_159 ),
	.F(\top/processor/sha_core/n3864_107 )
);
defparam \top/processor/sha_core/n3864_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3720_s138  (
	.I0(\top/processor/sha_core/n3622_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [16]),
	.I3(\top/processor/sha_core/w[12] [16]),
	.F(\top/processor/sha_core/n3622_155 )
);
defparam \top/processor/sha_core/n3720_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s138  (
	.I0(\top/processor/sha_core/n3623_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [15]),
	.I3(\top/processor/sha_core/w[12] [15]),
	.F(\top/processor/sha_core/n3623_155 )
);
defparam \top/processor/sha_core/n3721_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s138  (
	.I0(\top/processor/sha_core/n3624_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [14]),
	.I3(\top/processor/sha_core/w[12] [14]),
	.F(\top/processor/sha_core/n3624_155 )
);
defparam \top/processor/sha_core/n3722_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s138  (
	.I0(\top/processor/sha_core/n3625_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [13]),
	.I3(\top/processor/sha_core/w[12] [13]),
	.F(\top/processor/sha_core/n3625_155 )
);
defparam \top/processor/sha_core/n3723_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s138  (
	.I0(\top/processor/sha_core/n3626_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [12]),
	.I3(\top/processor/sha_core/w[12] [12]),
	.F(\top/processor/sha_core/n3626_155 )
);
defparam \top/processor/sha_core/n3724_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s138  (
	.I0(\top/processor/sha_core/n3627_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [11]),
	.I3(\top/processor/sha_core/w[12] [11]),
	.F(\top/processor/sha_core/n3627_155 )
);
defparam \top/processor/sha_core/n3725_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s138  (
	.I0(\top/processor/sha_core/n3628_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [10]),
	.I3(\top/processor/sha_core/w[12] [10]),
	.F(\top/processor/sha_core/n3628_155 )
);
defparam \top/processor/sha_core/n3726_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s138  (
	.I0(\top/processor/sha_core/n3629_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [9]),
	.I3(\top/processor/sha_core/w[12] [9]),
	.F(\top/processor/sha_core/n3629_155 )
);
defparam \top/processor/sha_core/n3727_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s138  (
	.I0(\top/processor/sha_core/n3630_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [8]),
	.I3(\top/processor/sha_core/w[12] [8]),
	.F(\top/processor/sha_core/n3630_155 )
);
defparam \top/processor/sha_core/n3728_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s138  (
	.I0(\top/processor/sha_core/n3631_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [7]),
	.I3(\top/processor/sha_core/w[12] [7]),
	.F(\top/processor/sha_core/n3631_155 )
);
defparam \top/processor/sha_core/n3729_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s138  (
	.I0(\top/processor/sha_core/n3632_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [6]),
	.I3(\top/processor/sha_core/w[12] [6]),
	.F(\top/processor/sha_core/n3632_155 )
);
defparam \top/processor/sha_core/n3730_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s138  (
	.I0(\top/processor/sha_core/n3633_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [5]),
	.I3(\top/processor/sha_core/w[12] [5]),
	.F(\top/processor/sha_core/n3633_155 )
);
defparam \top/processor/sha_core/n3731_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s138  (
	.I0(\top/processor/sha_core/n3634_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [4]),
	.I3(\top/processor/sha_core/w[12] [4]),
	.F(\top/processor/sha_core/n3634_155 )
);
defparam \top/processor/sha_core/n3732_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s138  (
	.I0(\top/processor/sha_core/n3635_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [3]),
	.I3(\top/processor/sha_core/w[12] [3]),
	.F(\top/processor/sha_core/n3635_155 )
);
defparam \top/processor/sha_core/n3733_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s138  (
	.I0(\top/processor/sha_core/n3636_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [2]),
	.I3(\top/processor/sha_core/w[12] [2]),
	.F(\top/processor/sha_core/n3636_155 )
);
defparam \top/processor/sha_core/n3734_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s138  (
	.I0(\top/processor/sha_core/n3637_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [1]),
	.I3(\top/processor/sha_core/w[12] [1]),
	.F(\top/processor/sha_core/n3637_155 )
);
defparam \top/processor/sha_core/n3735_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s138  (
	.I0(\top/processor/sha_core/n3638_175 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[14] [0]),
	.I3(\top/processor/sha_core/w[12] [0]),
	.F(\top/processor/sha_core/n3638_155 )
);
defparam \top/processor/sha_core/n3736_s138 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3492_s184  (
	.I0(\top/processor/sha_core/n3492_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_161 ),
	.I3(\top/processor/sha_core/n3492_162 ),
	.F(\top/processor/sha_core/n3492_141 )
);
defparam \top/processor/sha_core/n3492_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s136  (
	.I0(\top/processor/sha_core/n3864_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_125 ),
	.I3(\top/processor/sha_core/n3492_162 ),
	.F(\top/processor/sha_core/n3864_109 )
);
defparam \top/processor/sha_core/n3864_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3492_s185  (
	.I0(\top/processor/sha_core/n3492_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_164 ),
	.I3(\top/processor/sha_core/n3492_165 ),
	.F(\top/processor/sha_core/n3492_143 )
);
defparam \top/processor/sha_core/n3492_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s137  (
	.I0(\top/processor/sha_core/n3864_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_127 ),
	.I3(\top/processor/sha_core/n3492_165 ),
	.F(\top/processor/sha_core/n3864_111 )
);
defparam \top/processor/sha_core/n3864_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s139  (
	.I0(\top/processor/sha_core/n3607_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [31]),
	.I3(\top/processor/sha_core/w[16] [31]),
	.F(\top/processor/sha_core/n3607_157 )
);
defparam \top/processor/sha_core/n3705_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s139  (
	.I0(\top/processor/sha_core/n3608_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [30]),
	.I3(\top/processor/sha_core/w[16] [30]),
	.F(\top/processor/sha_core/n3608_157 )
);
defparam \top/processor/sha_core/n3706_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s139  (
	.I0(\top/processor/sha_core/n3609_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [29]),
	.I3(\top/processor/sha_core/w[16] [29]),
	.F(\top/processor/sha_core/n3609_157 )
);
defparam \top/processor/sha_core/n3707_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s139  (
	.I0(\top/processor/sha_core/n3610_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [28]),
	.I3(\top/processor/sha_core/w[16] [28]),
	.F(\top/processor/sha_core/n3610_157 )
);
defparam \top/processor/sha_core/n3708_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s139  (
	.I0(\top/processor/sha_core/n3611_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [27]),
	.I3(\top/processor/sha_core/w[16] [27]),
	.F(\top/processor/sha_core/n3611_157 )
);
defparam \top/processor/sha_core/n3709_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s139  (
	.I0(\top/processor/sha_core/n3612_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [26]),
	.I3(\top/processor/sha_core/w[16] [26]),
	.F(\top/processor/sha_core/n3612_157 )
);
defparam \top/processor/sha_core/n3710_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s139  (
	.I0(\top/processor/sha_core/n3613_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [25]),
	.I3(\top/processor/sha_core/w[16] [25]),
	.F(\top/processor/sha_core/n3613_157 )
);
defparam \top/processor/sha_core/n3711_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s139  (
	.I0(\top/processor/sha_core/n3614_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [24]),
	.I3(\top/processor/sha_core/w[16] [24]),
	.F(\top/processor/sha_core/n3614_157 )
);
defparam \top/processor/sha_core/n3712_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s139  (
	.I0(\top/processor/sha_core/n3615_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [23]),
	.I3(\top/processor/sha_core/w[16] [23]),
	.F(\top/processor/sha_core/n3615_157 )
);
defparam \top/processor/sha_core/n3713_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s139  (
	.I0(\top/processor/sha_core/n3616_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [22]),
	.I3(\top/processor/sha_core/w[16] [22]),
	.F(\top/processor/sha_core/n3616_157 )
);
defparam \top/processor/sha_core/n3714_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s139  (
	.I0(\top/processor/sha_core/n3617_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [21]),
	.I3(\top/processor/sha_core/w[16] [21]),
	.F(\top/processor/sha_core/n3617_157 )
);
defparam \top/processor/sha_core/n3715_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3492_s186  (
	.I0(\top/processor/sha_core/n3492_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_167 ),
	.I3(\top/processor/sha_core/n3492_168 ),
	.F(\top/processor/sha_core/n3492_145 )
);
defparam \top/processor/sha_core/n3492_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s138  (
	.I0(\top/processor/sha_core/n3864_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_129 ),
	.I3(\top/processor/sha_core/n3492_168 ),
	.F(\top/processor/sha_core/n3864_113 )
);
defparam \top/processor/sha_core/n3864_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3716_s139  (
	.I0(\top/processor/sha_core/n3618_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [20]),
	.I3(\top/processor/sha_core/w[16] [20]),
	.F(\top/processor/sha_core/n3618_157 )
);
defparam \top/processor/sha_core/n3716_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s139  (
	.I0(\top/processor/sha_core/n3619_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [19]),
	.I3(\top/processor/sha_core/w[16] [19]),
	.F(\top/processor/sha_core/n3619_157 )
);
defparam \top/processor/sha_core/n3717_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s139  (
	.I0(\top/processor/sha_core/n3620_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [18]),
	.I3(\top/processor/sha_core/w[16] [18]),
	.F(\top/processor/sha_core/n3620_157 )
);
defparam \top/processor/sha_core/n3718_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s139  (
	.I0(\top/processor/sha_core/n3621_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [17]),
	.I3(\top/processor/sha_core/w[16] [17]),
	.F(\top/processor/sha_core/n3621_157 )
);
defparam \top/processor/sha_core/n3719_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s139  (
	.I0(\top/processor/sha_core/n3622_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [16]),
	.I3(\top/processor/sha_core/w[16] [16]),
	.F(\top/processor/sha_core/n3622_157 )
);
defparam \top/processor/sha_core/n3720_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s139  (
	.I0(\top/processor/sha_core/n3623_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [15]),
	.I3(\top/processor/sha_core/w[16] [15]),
	.F(\top/processor/sha_core/n3623_157 )
);
defparam \top/processor/sha_core/n3721_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s139  (
	.I0(\top/processor/sha_core/n3624_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [14]),
	.I3(\top/processor/sha_core/w[16] [14]),
	.F(\top/processor/sha_core/n3624_157 )
);
defparam \top/processor/sha_core/n3722_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s139  (
	.I0(\top/processor/sha_core/n3625_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [13]),
	.I3(\top/processor/sha_core/w[16] [13]),
	.F(\top/processor/sha_core/n3625_157 )
);
defparam \top/processor/sha_core/n3723_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s139  (
	.I0(\top/processor/sha_core/n3626_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [12]),
	.I3(\top/processor/sha_core/w[16] [12]),
	.F(\top/processor/sha_core/n3626_157 )
);
defparam \top/processor/sha_core/n3724_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s139  (
	.I0(\top/processor/sha_core/n3627_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [11]),
	.I3(\top/processor/sha_core/w[16] [11]),
	.F(\top/processor/sha_core/n3627_157 )
);
defparam \top/processor/sha_core/n3725_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s139  (
	.I0(\top/processor/sha_core/n3628_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [10]),
	.I3(\top/processor/sha_core/w[16] [10]),
	.F(\top/processor/sha_core/n3628_157 )
);
defparam \top/processor/sha_core/n3726_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s139  (
	.I0(\top/processor/sha_core/n3629_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [9]),
	.I3(\top/processor/sha_core/w[16] [9]),
	.F(\top/processor/sha_core/n3629_157 )
);
defparam \top/processor/sha_core/n3727_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s139  (
	.I0(\top/processor/sha_core/n3630_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [8]),
	.I3(\top/processor/sha_core/w[16] [8]),
	.F(\top/processor/sha_core/n3630_157 )
);
defparam \top/processor/sha_core/n3728_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s139  (
	.I0(\top/processor/sha_core/n3631_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [7]),
	.I3(\top/processor/sha_core/w[16] [7]),
	.F(\top/processor/sha_core/n3631_157 )
);
defparam \top/processor/sha_core/n3729_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s139  (
	.I0(\top/processor/sha_core/n3632_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [6]),
	.I3(\top/processor/sha_core/w[16] [6]),
	.F(\top/processor/sha_core/n3632_157 )
);
defparam \top/processor/sha_core/n3730_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s139  (
	.I0(\top/processor/sha_core/n3633_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [5]),
	.I3(\top/processor/sha_core/w[16] [5]),
	.F(\top/processor/sha_core/n3633_157 )
);
defparam \top/processor/sha_core/n3731_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s139  (
	.I0(\top/processor/sha_core/n3634_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [4]),
	.I3(\top/processor/sha_core/w[16] [4]),
	.F(\top/processor/sha_core/n3634_157 )
);
defparam \top/processor/sha_core/n3732_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s139  (
	.I0(\top/processor/sha_core/n3635_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [3]),
	.I3(\top/processor/sha_core/w[16] [3]),
	.F(\top/processor/sha_core/n3635_157 )
);
defparam \top/processor/sha_core/n3733_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s139  (
	.I0(\top/processor/sha_core/n3636_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [2]),
	.I3(\top/processor/sha_core/w[16] [2]),
	.F(\top/processor/sha_core/n3636_157 )
);
defparam \top/processor/sha_core/n3734_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s139  (
	.I0(\top/processor/sha_core/n3637_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [1]),
	.I3(\top/processor/sha_core/w[16] [1]),
	.F(\top/processor/sha_core/n3637_157 )
);
defparam \top/processor/sha_core/n3735_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3492_s187  (
	.I0(\top/processor/sha_core/n3492_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_170 ),
	.I3(\top/processor/sha_core/n3492_171 ),
	.F(\top/processor/sha_core/n3492_147 )
);
defparam \top/processor/sha_core/n3492_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3864_s139  (
	.I0(\top/processor/sha_core/n3864_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3864_131 ),
	.I3(\top/processor/sha_core/n3492_171 ),
	.F(\top/processor/sha_core/n3864_115 )
);
defparam \top/processor/sha_core/n3864_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s183  (
	.I0(\top/processor/sha_core/n3488_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_167 ),
	.I3(\top/processor/sha_core/n3488_168 ),
	.F(\top/processor/sha_core/n3488_145 )
);
defparam \top/processor/sha_core/n3488_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s135  (
	.I0(\top/processor/sha_core/n3860_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_129 ),
	.I3(\top/processor/sha_core/n3488_168 ),
	.F(\top/processor/sha_core/n3860_113 )
);
defparam \top/processor/sha_core/n3860_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3736_s139  (
	.I0(\top/processor/sha_core/n3638_176 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[18] [0]),
	.I3(\top/processor/sha_core/w[16] [0]),
	.F(\top/processor/sha_core/n3638_157 )
);
defparam \top/processor/sha_core/n3736_s139 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s180  (
	.I0(\top/processor/sha_core/n3493_148 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_149 ),
	.I3(\top/processor/sha_core/n3493_150 ),
	.F(\top/processor/sha_core/n3493_133 )
);
defparam \top/processor/sha_core/n3493_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s132  (
	.I0(\top/processor/sha_core/n3865_116 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_117 ),
	.I3(\top/processor/sha_core/n3493_150 ),
	.F(\top/processor/sha_core/n3865_101 )
);
defparam \top/processor/sha_core/n3865_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s140  (
	.I0(\top/processor/sha_core/n3607_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [31]),
	.I3(\top/processor/sha_core/w[20] [31]),
	.F(\top/processor/sha_core/n3607_159 )
);
defparam \top/processor/sha_core/n3705_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s140  (
	.I0(\top/processor/sha_core/n3608_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [30]),
	.I3(\top/processor/sha_core/w[20] [30]),
	.F(\top/processor/sha_core/n3608_159 )
);
defparam \top/processor/sha_core/n3706_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s140  (
	.I0(\top/processor/sha_core/n3609_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [29]),
	.I3(\top/processor/sha_core/w[20] [29]),
	.F(\top/processor/sha_core/n3609_159 )
);
defparam \top/processor/sha_core/n3707_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s140  (
	.I0(\top/processor/sha_core/n3610_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [28]),
	.I3(\top/processor/sha_core/w[20] [28]),
	.F(\top/processor/sha_core/n3610_159 )
);
defparam \top/processor/sha_core/n3708_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s140  (
	.I0(\top/processor/sha_core/n3611_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [27]),
	.I3(\top/processor/sha_core/w[20] [27]),
	.F(\top/processor/sha_core/n3611_159 )
);
defparam \top/processor/sha_core/n3709_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s140  (
	.I0(\top/processor/sha_core/n3612_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [26]),
	.I3(\top/processor/sha_core/w[20] [26]),
	.F(\top/processor/sha_core/n3612_159 )
);
defparam \top/processor/sha_core/n3710_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s140  (
	.I0(\top/processor/sha_core/n3613_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [25]),
	.I3(\top/processor/sha_core/w[20] [25]),
	.F(\top/processor/sha_core/n3613_159 )
);
defparam \top/processor/sha_core/n3711_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s181  (
	.I0(\top/processor/sha_core/n3493_151 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_152 ),
	.I3(\top/processor/sha_core/n3493_153 ),
	.F(\top/processor/sha_core/n3493_135 )
);
defparam \top/processor/sha_core/n3493_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s133  (
	.I0(\top/processor/sha_core/n3865_118 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_119 ),
	.I3(\top/processor/sha_core/n3493_153 ),
	.F(\top/processor/sha_core/n3865_103 )
);
defparam \top/processor/sha_core/n3865_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3712_s140  (
	.I0(\top/processor/sha_core/n3614_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [24]),
	.I3(\top/processor/sha_core/w[20] [24]),
	.F(\top/processor/sha_core/n3614_159 )
);
defparam \top/processor/sha_core/n3712_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s140  (
	.I0(\top/processor/sha_core/n3615_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [23]),
	.I3(\top/processor/sha_core/w[20] [23]),
	.F(\top/processor/sha_core/n3615_159 )
);
defparam \top/processor/sha_core/n3713_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s140  (
	.I0(\top/processor/sha_core/n3616_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [22]),
	.I3(\top/processor/sha_core/w[20] [22]),
	.F(\top/processor/sha_core/n3616_159 )
);
defparam \top/processor/sha_core/n3714_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s140  (
	.I0(\top/processor/sha_core/n3617_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [21]),
	.I3(\top/processor/sha_core/w[20] [21]),
	.F(\top/processor/sha_core/n3617_159 )
);
defparam \top/processor/sha_core/n3715_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s140  (
	.I0(\top/processor/sha_core/n3618_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [20]),
	.I3(\top/processor/sha_core/w[20] [20]),
	.F(\top/processor/sha_core/n3618_159 )
);
defparam \top/processor/sha_core/n3716_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s140  (
	.I0(\top/processor/sha_core/n3619_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [19]),
	.I3(\top/processor/sha_core/w[20] [19]),
	.F(\top/processor/sha_core/n3619_159 )
);
defparam \top/processor/sha_core/n3717_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s140  (
	.I0(\top/processor/sha_core/n3620_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [18]),
	.I3(\top/processor/sha_core/w[20] [18]),
	.F(\top/processor/sha_core/n3620_159 )
);
defparam \top/processor/sha_core/n3718_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s140  (
	.I0(\top/processor/sha_core/n3621_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [17]),
	.I3(\top/processor/sha_core/w[20] [17]),
	.F(\top/processor/sha_core/n3621_159 )
);
defparam \top/processor/sha_core/n3719_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s140  (
	.I0(\top/processor/sha_core/n3622_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [16]),
	.I3(\top/processor/sha_core/w[20] [16]),
	.F(\top/processor/sha_core/n3622_159 )
);
defparam \top/processor/sha_core/n3720_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s140  (
	.I0(\top/processor/sha_core/n3623_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [15]),
	.I3(\top/processor/sha_core/w[20] [15]),
	.F(\top/processor/sha_core/n3623_159 )
);
defparam \top/processor/sha_core/n3721_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s140  (
	.I0(\top/processor/sha_core/n3624_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [14]),
	.I3(\top/processor/sha_core/w[20] [14]),
	.F(\top/processor/sha_core/n3624_159 )
);
defparam \top/processor/sha_core/n3722_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s140  (
	.I0(\top/processor/sha_core/n3625_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [13]),
	.I3(\top/processor/sha_core/w[20] [13]),
	.F(\top/processor/sha_core/n3625_159 )
);
defparam \top/processor/sha_core/n3723_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s140  (
	.I0(\top/processor/sha_core/n3626_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [12]),
	.I3(\top/processor/sha_core/w[20] [12]),
	.F(\top/processor/sha_core/n3626_159 )
);
defparam \top/processor/sha_core/n3724_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s140  (
	.I0(\top/processor/sha_core/n3627_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [11]),
	.I3(\top/processor/sha_core/w[20] [11]),
	.F(\top/processor/sha_core/n3627_159 )
);
defparam \top/processor/sha_core/n3725_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s140  (
	.I0(\top/processor/sha_core/n3628_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [10]),
	.I3(\top/processor/sha_core/w[20] [10]),
	.F(\top/processor/sha_core/n3628_159 )
);
defparam \top/processor/sha_core/n3726_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s140  (
	.I0(\top/processor/sha_core/n3629_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [9]),
	.I3(\top/processor/sha_core/w[20] [9]),
	.F(\top/processor/sha_core/n3629_159 )
);
defparam \top/processor/sha_core/n3727_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s140  (
	.I0(\top/processor/sha_core/n3630_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [8]),
	.I3(\top/processor/sha_core/w[20] [8]),
	.F(\top/processor/sha_core/n3630_159 )
);
defparam \top/processor/sha_core/n3728_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s140  (
	.I0(\top/processor/sha_core/n3631_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [7]),
	.I3(\top/processor/sha_core/w[20] [7]),
	.F(\top/processor/sha_core/n3631_159 )
);
defparam \top/processor/sha_core/n3729_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s140  (
	.I0(\top/processor/sha_core/n3632_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [6]),
	.I3(\top/processor/sha_core/w[20] [6]),
	.F(\top/processor/sha_core/n3632_159 )
);
defparam \top/processor/sha_core/n3730_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s140  (
	.I0(\top/processor/sha_core/n3633_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [5]),
	.I3(\top/processor/sha_core/w[20] [5]),
	.F(\top/processor/sha_core/n3633_159 )
);
defparam \top/processor/sha_core/n3731_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s182  (
	.I0(\top/processor/sha_core/n3493_154 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_155 ),
	.I3(\top/processor/sha_core/n3493_156 ),
	.F(\top/processor/sha_core/n3493_137 )
);
defparam \top/processor/sha_core/n3493_s182 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s134  (
	.I0(\top/processor/sha_core/n3865_120 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_121 ),
	.I3(\top/processor/sha_core/n3493_156 ),
	.F(\top/processor/sha_core/n3865_105 )
);
defparam \top/processor/sha_core/n3865_s134 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3732_s140  (
	.I0(\top/processor/sha_core/n3634_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [4]),
	.I3(\top/processor/sha_core/w[20] [4]),
	.F(\top/processor/sha_core/n3634_159 )
);
defparam \top/processor/sha_core/n3732_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s140  (
	.I0(\top/processor/sha_core/n3635_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [3]),
	.I3(\top/processor/sha_core/w[20] [3]),
	.F(\top/processor/sha_core/n3635_159 )
);
defparam \top/processor/sha_core/n3733_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s140  (
	.I0(\top/processor/sha_core/n3636_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [2]),
	.I3(\top/processor/sha_core/w[20] [2]),
	.F(\top/processor/sha_core/n3636_159 )
);
defparam \top/processor/sha_core/n3734_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s140  (
	.I0(\top/processor/sha_core/n3637_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [1]),
	.I3(\top/processor/sha_core/w[20] [1]),
	.F(\top/processor/sha_core/n3637_159 )
);
defparam \top/processor/sha_core/n3735_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s140  (
	.I0(\top/processor/sha_core/n3638_177 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[22] [0]),
	.I3(\top/processor/sha_core/w[20] [0]),
	.F(\top/processor/sha_core/n3638_159 )
);
defparam \top/processor/sha_core/n3736_s140 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s183  (
	.I0(\top/processor/sha_core/n3493_157 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_158 ),
	.I3(\top/processor/sha_core/n3493_159 ),
	.F(\top/processor/sha_core/n3493_139 )
);
defparam \top/processor/sha_core/n3493_s183 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s135  (
	.I0(\top/processor/sha_core/n3865_122 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_123 ),
	.I3(\top/processor/sha_core/n3493_159 ),
	.F(\top/processor/sha_core/n3865_107 )
);
defparam \top/processor/sha_core/n3865_s135 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s141  (
	.I0(\top/processor/sha_core/n3607_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [31]),
	.I3(\top/processor/sha_core/w[24] [31]),
	.F(\top/processor/sha_core/n3607_161 )
);
defparam \top/processor/sha_core/n3705_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s141  (
	.I0(\top/processor/sha_core/n3608_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [30]),
	.I3(\top/processor/sha_core/w[24] [30]),
	.F(\top/processor/sha_core/n3608_161 )
);
defparam \top/processor/sha_core/n3706_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s141  (
	.I0(\top/processor/sha_core/n3609_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [29]),
	.I3(\top/processor/sha_core/w[24] [29]),
	.F(\top/processor/sha_core/n3609_161 )
);
defparam \top/processor/sha_core/n3707_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s184  (
	.I0(\top/processor/sha_core/n3493_160 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_161 ),
	.I3(\top/processor/sha_core/n3493_162 ),
	.F(\top/processor/sha_core/n3493_141 )
);
defparam \top/processor/sha_core/n3493_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s136  (
	.I0(\top/processor/sha_core/n3865_124 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_125 ),
	.I3(\top/processor/sha_core/n3493_162 ),
	.F(\top/processor/sha_core/n3865_109 )
);
defparam \top/processor/sha_core/n3865_s136 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3708_s141  (
	.I0(\top/processor/sha_core/n3610_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [28]),
	.I3(\top/processor/sha_core/w[24] [28]),
	.F(\top/processor/sha_core/n3610_161 )
);
defparam \top/processor/sha_core/n3708_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s141  (
	.I0(\top/processor/sha_core/n3611_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [27]),
	.I3(\top/processor/sha_core/w[24] [27]),
	.F(\top/processor/sha_core/n3611_161 )
);
defparam \top/processor/sha_core/n3709_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s141  (
	.I0(\top/processor/sha_core/n3612_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [26]),
	.I3(\top/processor/sha_core/w[24] [26]),
	.F(\top/processor/sha_core/n3612_161 )
);
defparam \top/processor/sha_core/n3710_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s141  (
	.I0(\top/processor/sha_core/n3613_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [25]),
	.I3(\top/processor/sha_core/w[24] [25]),
	.F(\top/processor/sha_core/n3613_161 )
);
defparam \top/processor/sha_core/n3711_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s141  (
	.I0(\top/processor/sha_core/n3614_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [24]),
	.I3(\top/processor/sha_core/w[24] [24]),
	.F(\top/processor/sha_core/n3614_161 )
);
defparam \top/processor/sha_core/n3712_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s141  (
	.I0(\top/processor/sha_core/n3615_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [23]),
	.I3(\top/processor/sha_core/w[24] [23]),
	.F(\top/processor/sha_core/n3615_161 )
);
defparam \top/processor/sha_core/n3713_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s141  (
	.I0(\top/processor/sha_core/n3616_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [22]),
	.I3(\top/processor/sha_core/w[24] [22]),
	.F(\top/processor/sha_core/n3616_161 )
);
defparam \top/processor/sha_core/n3714_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s141  (
	.I0(\top/processor/sha_core/n3617_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [21]),
	.I3(\top/processor/sha_core/w[24] [21]),
	.F(\top/processor/sha_core/n3617_161 )
);
defparam \top/processor/sha_core/n3715_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s141  (
	.I0(\top/processor/sha_core/n3618_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [20]),
	.I3(\top/processor/sha_core/w[24] [20]),
	.F(\top/processor/sha_core/n3618_161 )
);
defparam \top/processor/sha_core/n3716_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s141  (
	.I0(\top/processor/sha_core/n3619_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [19]),
	.I3(\top/processor/sha_core/w[24] [19]),
	.F(\top/processor/sha_core/n3619_161 )
);
defparam \top/processor/sha_core/n3717_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s141  (
	.I0(\top/processor/sha_core/n3620_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [18]),
	.I3(\top/processor/sha_core/w[24] [18]),
	.F(\top/processor/sha_core/n3620_161 )
);
defparam \top/processor/sha_core/n3718_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s141  (
	.I0(\top/processor/sha_core/n3621_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [17]),
	.I3(\top/processor/sha_core/w[24] [17]),
	.F(\top/processor/sha_core/n3621_161 )
);
defparam \top/processor/sha_core/n3719_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s141  (
	.I0(\top/processor/sha_core/n3622_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [16]),
	.I3(\top/processor/sha_core/w[24] [16]),
	.F(\top/processor/sha_core/n3622_161 )
);
defparam \top/processor/sha_core/n3720_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s141  (
	.I0(\top/processor/sha_core/n3623_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [15]),
	.I3(\top/processor/sha_core/w[24] [15]),
	.F(\top/processor/sha_core/n3623_161 )
);
defparam \top/processor/sha_core/n3721_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s141  (
	.I0(\top/processor/sha_core/n3624_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [14]),
	.I3(\top/processor/sha_core/w[24] [14]),
	.F(\top/processor/sha_core/n3624_161 )
);
defparam \top/processor/sha_core/n3722_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s141  (
	.I0(\top/processor/sha_core/n3625_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [13]),
	.I3(\top/processor/sha_core/w[24] [13]),
	.F(\top/processor/sha_core/n3625_161 )
);
defparam \top/processor/sha_core/n3723_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3724_s141  (
	.I0(\top/processor/sha_core/n3626_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [12]),
	.I3(\top/processor/sha_core/w[24] [12]),
	.F(\top/processor/sha_core/n3626_161 )
);
defparam \top/processor/sha_core/n3724_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s141  (
	.I0(\top/processor/sha_core/n3627_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [11]),
	.I3(\top/processor/sha_core/w[24] [11]),
	.F(\top/processor/sha_core/n3627_161 )
);
defparam \top/processor/sha_core/n3725_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s141  (
	.I0(\top/processor/sha_core/n3628_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [10]),
	.I3(\top/processor/sha_core/w[24] [10]),
	.F(\top/processor/sha_core/n3628_161 )
);
defparam \top/processor/sha_core/n3726_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s141  (
	.I0(\top/processor/sha_core/n3629_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [9]),
	.I3(\top/processor/sha_core/w[24] [9]),
	.F(\top/processor/sha_core/n3629_161 )
);
defparam \top/processor/sha_core/n3727_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s185  (
	.I0(\top/processor/sha_core/n3493_163 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_164 ),
	.I3(\top/processor/sha_core/n3493_165 ),
	.F(\top/processor/sha_core/n3493_143 )
);
defparam \top/processor/sha_core/n3493_s185 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s137  (
	.I0(\top/processor/sha_core/n3865_126 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_127 ),
	.I3(\top/processor/sha_core/n3493_165 ),
	.F(\top/processor/sha_core/n3865_111 )
);
defparam \top/processor/sha_core/n3865_s137 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3728_s141  (
	.I0(\top/processor/sha_core/n3630_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [8]),
	.I3(\top/processor/sha_core/w[24] [8]),
	.F(\top/processor/sha_core/n3630_161 )
);
defparam \top/processor/sha_core/n3728_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s141  (
	.I0(\top/processor/sha_core/n3631_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [7]),
	.I3(\top/processor/sha_core/w[24] [7]),
	.F(\top/processor/sha_core/n3631_161 )
);
defparam \top/processor/sha_core/n3729_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s141  (
	.I0(\top/processor/sha_core/n3632_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [6]),
	.I3(\top/processor/sha_core/w[24] [6]),
	.F(\top/processor/sha_core/n3632_161 )
);
defparam \top/processor/sha_core/n3730_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s141  (
	.I0(\top/processor/sha_core/n3633_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [5]),
	.I3(\top/processor/sha_core/w[24] [5]),
	.F(\top/processor/sha_core/n3633_161 )
);
defparam \top/processor/sha_core/n3731_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s141  (
	.I0(\top/processor/sha_core/n3634_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [4]),
	.I3(\top/processor/sha_core/w[24] [4]),
	.F(\top/processor/sha_core/n3634_161 )
);
defparam \top/processor/sha_core/n3732_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s141  (
	.I0(\top/processor/sha_core/n3635_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [3]),
	.I3(\top/processor/sha_core/w[24] [3]),
	.F(\top/processor/sha_core/n3635_161 )
);
defparam \top/processor/sha_core/n3733_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s141  (
	.I0(\top/processor/sha_core/n3636_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [2]),
	.I3(\top/processor/sha_core/w[24] [2]),
	.F(\top/processor/sha_core/n3636_161 )
);
defparam \top/processor/sha_core/n3734_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s141  (
	.I0(\top/processor/sha_core/n3637_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [1]),
	.I3(\top/processor/sha_core/w[24] [1]),
	.F(\top/processor/sha_core/n3637_161 )
);
defparam \top/processor/sha_core/n3735_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s141  (
	.I0(\top/processor/sha_core/n3638_178 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[26] [0]),
	.I3(\top/processor/sha_core/w[24] [0]),
	.F(\top/processor/sha_core/n3638_161 )
);
defparam \top/processor/sha_core/n3736_s141 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3493_s186  (
	.I0(\top/processor/sha_core/n3493_166 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_167 ),
	.I3(\top/processor/sha_core/n3493_168 ),
	.F(\top/processor/sha_core/n3493_145 )
);
defparam \top/processor/sha_core/n3493_s186 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s138  (
	.I0(\top/processor/sha_core/n3865_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_129 ),
	.I3(\top/processor/sha_core/n3493_168 ),
	.F(\top/processor/sha_core/n3865_113 )
);
defparam \top/processor/sha_core/n3865_s138 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3493_s187  (
	.I0(\top/processor/sha_core/n3493_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_170 ),
	.I3(\top/processor/sha_core/n3493_171 ),
	.F(\top/processor/sha_core/n3493_147 )
);
defparam \top/processor/sha_core/n3493_s187 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3865_s139  (
	.I0(\top/processor/sha_core/n3865_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3865_131 ),
	.I3(\top/processor/sha_core/n3493_171 ),
	.F(\top/processor/sha_core/n3865_115 )
);
defparam \top/processor/sha_core/n3865_s139 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3705_s142  (
	.I0(\top/processor/sha_core/n3607_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [31]),
	.I3(\top/processor/sha_core/w[28] [31]),
	.F(\top/processor/sha_core/n3607_163 )
);
defparam \top/processor/sha_core/n3705_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3706_s142  (
	.I0(\top/processor/sha_core/n3608_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [30]),
	.I3(\top/processor/sha_core/w[28] [30]),
	.F(\top/processor/sha_core/n3608_163 )
);
defparam \top/processor/sha_core/n3706_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3707_s142  (
	.I0(\top/processor/sha_core/n3609_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [29]),
	.I3(\top/processor/sha_core/w[28] [29]),
	.F(\top/processor/sha_core/n3609_163 )
);
defparam \top/processor/sha_core/n3707_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3708_s142  (
	.I0(\top/processor/sha_core/n3610_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [28]),
	.I3(\top/processor/sha_core/w[28] [28]),
	.F(\top/processor/sha_core/n3610_163 )
);
defparam \top/processor/sha_core/n3708_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3709_s142  (
	.I0(\top/processor/sha_core/n3611_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [27]),
	.I3(\top/processor/sha_core/w[28] [27]),
	.F(\top/processor/sha_core/n3611_163 )
);
defparam \top/processor/sha_core/n3709_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3710_s142  (
	.I0(\top/processor/sha_core/n3612_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [26]),
	.I3(\top/processor/sha_core/w[28] [26]),
	.F(\top/processor/sha_core/n3612_163 )
);
defparam \top/processor/sha_core/n3710_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3711_s142  (
	.I0(\top/processor/sha_core/n3613_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [25]),
	.I3(\top/processor/sha_core/w[28] [25]),
	.F(\top/processor/sha_core/n3613_163 )
);
defparam \top/processor/sha_core/n3711_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3712_s142  (
	.I0(\top/processor/sha_core/n3614_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [24]),
	.I3(\top/processor/sha_core/w[28] [24]),
	.F(\top/processor/sha_core/n3614_163 )
);
defparam \top/processor/sha_core/n3712_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3713_s142  (
	.I0(\top/processor/sha_core/n3615_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [23]),
	.I3(\top/processor/sha_core/w[28] [23]),
	.F(\top/processor/sha_core/n3615_163 )
);
defparam \top/processor/sha_core/n3713_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3714_s142  (
	.I0(\top/processor/sha_core/n3616_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [22]),
	.I3(\top/processor/sha_core/w[28] [22]),
	.F(\top/processor/sha_core/n3616_163 )
);
defparam \top/processor/sha_core/n3714_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3715_s142  (
	.I0(\top/processor/sha_core/n3617_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [21]),
	.I3(\top/processor/sha_core/w[28] [21]),
	.F(\top/processor/sha_core/n3617_163 )
);
defparam \top/processor/sha_core/n3715_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3716_s142  (
	.I0(\top/processor/sha_core/n3618_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [20]),
	.I3(\top/processor/sha_core/w[28] [20]),
	.F(\top/processor/sha_core/n3618_163 )
);
defparam \top/processor/sha_core/n3716_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3717_s142  (
	.I0(\top/processor/sha_core/n3619_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [19]),
	.I3(\top/processor/sha_core/w[28] [19]),
	.F(\top/processor/sha_core/n3619_163 )
);
defparam \top/processor/sha_core/n3717_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3718_s142  (
	.I0(\top/processor/sha_core/n3620_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [18]),
	.I3(\top/processor/sha_core/w[28] [18]),
	.F(\top/processor/sha_core/n3620_163 )
);
defparam \top/processor/sha_core/n3718_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3719_s142  (
	.I0(\top/processor/sha_core/n3621_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [17]),
	.I3(\top/processor/sha_core/w[28] [17]),
	.F(\top/processor/sha_core/n3621_163 )
);
defparam \top/processor/sha_core/n3719_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3720_s142  (
	.I0(\top/processor/sha_core/n3622_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [16]),
	.I3(\top/processor/sha_core/w[28] [16]),
	.F(\top/processor/sha_core/n3622_163 )
);
defparam \top/processor/sha_core/n3720_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3721_s142  (
	.I0(\top/processor/sha_core/n3623_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [15]),
	.I3(\top/processor/sha_core/w[28] [15]),
	.F(\top/processor/sha_core/n3623_163 )
);
defparam \top/processor/sha_core/n3721_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3722_s142  (
	.I0(\top/processor/sha_core/n3624_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [14]),
	.I3(\top/processor/sha_core/w[28] [14]),
	.F(\top/processor/sha_core/n3624_163 )
);
defparam \top/processor/sha_core/n3722_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3723_s142  (
	.I0(\top/processor/sha_core/n3625_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [13]),
	.I3(\top/processor/sha_core/w[28] [13]),
	.F(\top/processor/sha_core/n3625_163 )
);
defparam \top/processor/sha_core/n3723_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s180  (
	.I0(\top/processor/sha_core/n3494_167 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_168 ),
	.I3(\top/processor/sha_core/n3494_169 ),
	.F(\top/processor/sha_core/n3494_145 )
);
defparam \top/processor/sha_core/n3494_s180 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s132  (
	.I0(\top/processor/sha_core/n3866_128 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_129 ),
	.I3(\top/processor/sha_core/n3494_169 ),
	.F(\top/processor/sha_core/n3866_113 )
);
defparam \top/processor/sha_core/n3866_s132 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3724_s142  (
	.I0(\top/processor/sha_core/n3626_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [12]),
	.I3(\top/processor/sha_core/w[28] [12]),
	.F(\top/processor/sha_core/n3626_163 )
);
defparam \top/processor/sha_core/n3724_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3725_s142  (
	.I0(\top/processor/sha_core/n3627_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [11]),
	.I3(\top/processor/sha_core/w[28] [11]),
	.F(\top/processor/sha_core/n3627_163 )
);
defparam \top/processor/sha_core/n3725_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3726_s142  (
	.I0(\top/processor/sha_core/n3628_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [10]),
	.I3(\top/processor/sha_core/w[28] [10]),
	.F(\top/processor/sha_core/n3628_163 )
);
defparam \top/processor/sha_core/n3726_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3727_s142  (
	.I0(\top/processor/sha_core/n3629_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [9]),
	.I3(\top/processor/sha_core/w[28] [9]),
	.F(\top/processor/sha_core/n3629_163 )
);
defparam \top/processor/sha_core/n3727_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3728_s142  (
	.I0(\top/processor/sha_core/n3630_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [8]),
	.I3(\top/processor/sha_core/w[28] [8]),
	.F(\top/processor/sha_core/n3630_163 )
);
defparam \top/processor/sha_core/n3728_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3729_s142  (
	.I0(\top/processor/sha_core/n3631_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [7]),
	.I3(\top/processor/sha_core/w[28] [7]),
	.F(\top/processor/sha_core/n3631_163 )
);
defparam \top/processor/sha_core/n3729_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3730_s142  (
	.I0(\top/processor/sha_core/n3632_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [6]),
	.I3(\top/processor/sha_core/w[28] [6]),
	.F(\top/processor/sha_core/n3632_163 )
);
defparam \top/processor/sha_core/n3730_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3731_s142  (
	.I0(\top/processor/sha_core/n3633_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [5]),
	.I3(\top/processor/sha_core/w[28] [5]),
	.F(\top/processor/sha_core/n3633_163 )
);
defparam \top/processor/sha_core/n3731_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3732_s142  (
	.I0(\top/processor/sha_core/n3634_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [4]),
	.I3(\top/processor/sha_core/w[28] [4]),
	.F(\top/processor/sha_core/n3634_163 )
);
defparam \top/processor/sha_core/n3732_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3733_s142  (
	.I0(\top/processor/sha_core/n3635_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [3]),
	.I3(\top/processor/sha_core/w[28] [3]),
	.F(\top/processor/sha_core/n3635_163 )
);
defparam \top/processor/sha_core/n3733_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3734_s142  (
	.I0(\top/processor/sha_core/n3636_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [2]),
	.I3(\top/processor/sha_core/w[28] [2]),
	.F(\top/processor/sha_core/n3636_163 )
);
defparam \top/processor/sha_core/n3734_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3735_s142  (
	.I0(\top/processor/sha_core/n3637_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [1]),
	.I3(\top/processor/sha_core/w[28] [1]),
	.F(\top/processor/sha_core/n3637_163 )
);
defparam \top/processor/sha_core/n3735_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3736_s142  (
	.I0(\top/processor/sha_core/n3638_179 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[30] [0]),
	.I3(\top/processor/sha_core/w[28] [0]),
	.F(\top/processor/sha_core/n3638_163 )
);
defparam \top/processor/sha_core/n3736_s142 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s181  (
	.I0(\top/processor/sha_core/n3494_170 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_171 ),
	.I3(\top/processor/sha_core/n3494_172 ),
	.F(\top/processor/sha_core/n3494_147 )
);
defparam \top/processor/sha_core/n3494_s181 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3866_s133  (
	.I0(\top/processor/sha_core/n3866_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3866_131 ),
	.I3(\top/processor/sha_core/n3494_172 ),
	.F(\top/processor/sha_core/n3866_115 )
);
defparam \top/processor/sha_core/n3866_s133 .INIT=16'hE6A2;
LUT4 \top/processor/sha_core/n3488_s184  (
	.I0(\top/processor/sha_core/n3488_169 ),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_170 ),
	.I3(\top/processor/sha_core/n3488_171 ),
	.F(\top/processor/sha_core/n3488_147 )
);
defparam \top/processor/sha_core/n3488_s184 .INIT=16'hEA62;
LUT4 \top/processor/sha_core/n3860_s136  (
	.I0(\top/processor/sha_core/n3860_130 ),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/n3860_131 ),
	.I3(\top/processor/sha_core/n3488_171 ),
	.F(\top/processor/sha_core/n3860_115 )
);
defparam \top/processor/sha_core/n3860_s136 .INIT=16'hD591;
LUT4 \top/processor/sha_core/n3494_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_117 ),
	.I3(\top/processor/sha_core/n3494_173 ),
	.F(\top/processor/sha_core/n3494_149 )
);
defparam \top/processor/sha_core/n3494_s135 .INIT=16'h7362;
LUT3 \top/processor/sha_core/n3494_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [25]),
	.I2(\top/processor/sha_core/w[17] [25]),
	.F(\top/processor/sha_core/n3494_150 )
);
defparam \top/processor/sha_core/n3494_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [25]),
	.I2(\top/processor/sha_core/w[21] [25]),
	.F(\top/processor/sha_core/n3494_151 )
);
defparam \top/processor/sha_core/n3494_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_173 ),
	.I3(\top/processor/sha_core/n3494_150 ),
	.F(\top/processor/sha_core/n3866_116 )
);
defparam \top/processor/sha_core/n3866_s103 .INIT=16'h7362;
LUT3 \top/processor/sha_core/n3866_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [25]),
	.I2(\top/processor/sha_core/w[23] [25]),
	.F(\top/processor/sha_core/n3866_117 )
);
defparam \top/processor/sha_core/n3866_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s143  (
	.I0(\top/processor/sha_core/n3453_7 ),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/w[32] [31]),
	.I3(\top/processor/sha_core/w[33] [31]),
	.F(\top/processor/sha_core/n3607_164 )
);
defparam \top/processor/sha_core/n3607_s143 .INIT=16'h2637;
LUT4 \top/processor/sha_core/n3608_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [30]),
	.I3(\top/processor/sha_core/w[33] [30]),
	.F(\top/processor/sha_core/n3608_164 )
);
defparam \top/processor/sha_core/n3608_s143 .INIT=16'h2637;
LUT4 \top/processor/sha_core/n3609_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [29]),
	.I3(\top/processor/sha_core/w[33] [29]),
	.F(\top/processor/sha_core/n3609_164 )
);
defparam \top/processor/sha_core/n3609_s143 .INIT=16'h2637;
LUT4 \top/processor/sha_core/n3610_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [28]),
	.I3(\top/processor/sha_core/w[33] [28]),
	.F(\top/processor/sha_core/n3610_164 )
);
defparam \top/processor/sha_core/n3610_s143 .INIT=16'h2637;
LUT4 \top/processor/sha_core/n3611_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [27]),
	.I3(\top/processor/sha_core/w[33] [27]),
	.F(\top/processor/sha_core/n3611_164 )
);
defparam \top/processor/sha_core/n3611_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [26]),
	.I3(\top/processor/sha_core/w[33] [26]),
	.F(\top/processor/sha_core/n3612_164 )
);
defparam \top/processor/sha_core/n3612_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [25]),
	.I3(\top/processor/sha_core/w[33] [25]),
	.F(\top/processor/sha_core/n3613_164 )
);
defparam \top/processor/sha_core/n3613_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [24]),
	.I3(\top/processor/sha_core/w[33] [24]),
	.F(\top/processor/sha_core/n3614_164 )
);
defparam \top/processor/sha_core/n3614_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [23]),
	.I3(\top/processor/sha_core/w[33] [23]),
	.F(\top/processor/sha_core/n3615_164 )
);
defparam \top/processor/sha_core/n3615_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [22]),
	.I3(\top/processor/sha_core/w[33] [22]),
	.F(\top/processor/sha_core/n3616_164 )
);
defparam \top/processor/sha_core/n3616_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [21]),
	.I3(\top/processor/sha_core/w[33] [21]),
	.F(\top/processor/sha_core/n3617_164 )
);
defparam \top/processor/sha_core/n3617_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [20]),
	.I3(\top/processor/sha_core/w[33] [20]),
	.F(\top/processor/sha_core/n3618_164 )
);
defparam \top/processor/sha_core/n3618_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [19]),
	.I3(\top/processor/sha_core/w[33] [19]),
	.F(\top/processor/sha_core/n3619_164 )
);
defparam \top/processor/sha_core/n3619_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [18]),
	.I3(\top/processor/sha_core/w[33] [18]),
	.F(\top/processor/sha_core/n3620_164 )
);
defparam \top/processor/sha_core/n3620_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [17]),
	.I3(\top/processor/sha_core/w[33] [17]),
	.F(\top/processor/sha_core/n3621_164 )
);
defparam \top/processor/sha_core/n3621_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3494_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_119 ),
	.I3(\top/processor/sha_core/n3494_174 ),
	.F(\top/processor/sha_core/n3494_152 )
);
defparam \top/processor/sha_core/n3494_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [25]),
	.I2(\top/processor/sha_core/w[25] [25]),
	.F(\top/processor/sha_core/n3494_153 )
);
defparam \top/processor/sha_core/n3494_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [25]),
	.I2(\top/processor/sha_core/w[29] [25]),
	.F(\top/processor/sha_core/n3494_154 )
);
defparam \top/processor/sha_core/n3494_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_174 ),
	.I3(\top/processor/sha_core/n3494_153 ),
	.F(\top/processor/sha_core/n3866_118 )
);
defparam \top/processor/sha_core/n3866_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [25]),
	.I2(\top/processor/sha_core/w[31] [25]),
	.F(\top/processor/sha_core/n3866_119 )
);
defparam \top/processor/sha_core/n3866_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3622_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [16]),
	.I3(\top/processor/sha_core/w[33] [16]),
	.F(\top/processor/sha_core/n3622_164 )
);
defparam \top/processor/sha_core/n3622_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [15]),
	.I3(\top/processor/sha_core/w[33] [15]),
	.F(\top/processor/sha_core/n3623_164 )
);
defparam \top/processor/sha_core/n3623_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [14]),
	.I3(\top/processor/sha_core/w[33] [14]),
	.F(\top/processor/sha_core/n3624_164 )
);
defparam \top/processor/sha_core/n3624_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [13]),
	.I3(\top/processor/sha_core/w[33] [13]),
	.F(\top/processor/sha_core/n3625_164 )
);
defparam \top/processor/sha_core/n3625_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [12]),
	.I3(\top/processor/sha_core/w[33] [12]),
	.F(\top/processor/sha_core/n3626_164 )
);
defparam \top/processor/sha_core/n3626_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [11]),
	.I3(\top/processor/sha_core/w[33] [11]),
	.F(\top/processor/sha_core/n3627_164 )
);
defparam \top/processor/sha_core/n3627_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [10]),
	.I3(\top/processor/sha_core/w[33] [10]),
	.F(\top/processor/sha_core/n3628_164 )
);
defparam \top/processor/sha_core/n3628_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [9]),
	.I3(\top/processor/sha_core/w[33] [9]),
	.F(\top/processor/sha_core/n3629_164 )
);
defparam \top/processor/sha_core/n3629_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [8]),
	.I3(\top/processor/sha_core/w[33] [8]),
	.F(\top/processor/sha_core/n3630_164 )
);
defparam \top/processor/sha_core/n3630_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [7]),
	.I3(\top/processor/sha_core/w[33] [7]),
	.F(\top/processor/sha_core/n3631_164 )
);
defparam \top/processor/sha_core/n3631_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [6]),
	.I3(\top/processor/sha_core/w[33] [6]),
	.F(\top/processor/sha_core/n3632_164 )
);
defparam \top/processor/sha_core/n3632_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [5]),
	.I3(\top/processor/sha_core/w[33] [5]),
	.F(\top/processor/sha_core/n3633_164 )
);
defparam \top/processor/sha_core/n3633_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [4]),
	.I3(\top/processor/sha_core/w[33] [4]),
	.F(\top/processor/sha_core/n3634_164 )
);
defparam \top/processor/sha_core/n3634_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [3]),
	.I3(\top/processor/sha_core/w[33] [3]),
	.F(\top/processor/sha_core/n3635_164 )
);
defparam \top/processor/sha_core/n3635_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [2]),
	.I3(\top/processor/sha_core/w[33] [2]),
	.F(\top/processor/sha_core/n3636_164 )
);
defparam \top/processor/sha_core/n3636_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [1]),
	.I3(\top/processor/sha_core/w[33] [1]),
	.F(\top/processor/sha_core/n3637_164 )
);
defparam \top/processor/sha_core/n3637_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[35] [0]),
	.I3(\top/processor/sha_core/w[33] [0]),
	.F(\top/processor/sha_core/n3638_164 )
);
defparam \top/processor/sha_core/n3638_s143 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3494_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_121 ),
	.I3(\top/processor/sha_core/n3494_175 ),
	.F(\top/processor/sha_core/n3494_155 )
);
defparam \top/processor/sha_core/n3494_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [25]),
	.I2(\top/processor/sha_core/w[33] [25]),
	.F(\top/processor/sha_core/n3494_156 )
);
defparam \top/processor/sha_core/n3494_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [25]),
	.I2(\top/processor/sha_core/w[37] [25]),
	.F(\top/processor/sha_core/n3494_157 )
);
defparam \top/processor/sha_core/n3494_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_175 ),
	.I3(\top/processor/sha_core/n3494_156 ),
	.F(\top/processor/sha_core/n3866_120 )
);
defparam \top/processor/sha_core/n3866_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [25]),
	.I2(\top/processor/sha_core/w[39] [25]),
	.F(\top/processor/sha_core/n3866_121 )
);
defparam \top/processor/sha_core/n3866_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3494_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_123 ),
	.I3(\top/processor/sha_core/n3494_176 ),
	.F(\top/processor/sha_core/n3494_158 )
);
defparam \top/processor/sha_core/n3494_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [25]),
	.I2(\top/processor/sha_core/w[41] [25]),
	.F(\top/processor/sha_core/n3494_159 )
);
defparam \top/processor/sha_core/n3494_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [25]),
	.I2(\top/processor/sha_core/w[45] [25]),
	.F(\top/processor/sha_core/n3494_160 )
);
defparam \top/processor/sha_core/n3494_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_176 ),
	.I3(\top/processor/sha_core/n3494_159 ),
	.F(\top/processor/sha_core/n3866_122 )
);
defparam \top/processor/sha_core/n3866_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [25]),
	.I2(\top/processor/sha_core/w[47] [25]),
	.F(\top/processor/sha_core/n3866_123 )
);
defparam \top/processor/sha_core/n3866_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [31]),
	.I3(\top/processor/sha_core/w[37] [31]),
	.F(\top/processor/sha_core/n3607_165 )
);
defparam \top/processor/sha_core/n3607_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [30]),
	.I3(\top/processor/sha_core/w[37] [30]),
	.F(\top/processor/sha_core/n3608_165 )
);
defparam \top/processor/sha_core/n3608_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [29]),
	.I3(\top/processor/sha_core/w[37] [29]),
	.F(\top/processor/sha_core/n3609_165 )
);
defparam \top/processor/sha_core/n3609_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [28]),
	.I3(\top/processor/sha_core/w[37] [28]),
	.F(\top/processor/sha_core/n3610_165 )
);
defparam \top/processor/sha_core/n3610_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [27]),
	.I3(\top/processor/sha_core/w[37] [27]),
	.F(\top/processor/sha_core/n3611_165 )
);
defparam \top/processor/sha_core/n3611_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [26]),
	.I3(\top/processor/sha_core/w[37] [26]),
	.F(\top/processor/sha_core/n3612_165 )
);
defparam \top/processor/sha_core/n3612_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [25]),
	.I3(\top/processor/sha_core/w[37] [25]),
	.F(\top/processor/sha_core/n3613_165 )
);
defparam \top/processor/sha_core/n3613_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [24]),
	.I3(\top/processor/sha_core/w[37] [24]),
	.F(\top/processor/sha_core/n3614_165 )
);
defparam \top/processor/sha_core/n3614_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [23]),
	.I3(\top/processor/sha_core/w[37] [23]),
	.F(\top/processor/sha_core/n3615_165 )
);
defparam \top/processor/sha_core/n3615_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [22]),
	.I3(\top/processor/sha_core/w[37] [22]),
	.F(\top/processor/sha_core/n3616_165 )
);
defparam \top/processor/sha_core/n3616_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [21]),
	.I3(\top/processor/sha_core/w[37] [21]),
	.F(\top/processor/sha_core/n3617_165 )
);
defparam \top/processor/sha_core/n3617_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3494_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_125 ),
	.I3(\top/processor/sha_core/n3494_177 ),
	.F(\top/processor/sha_core/n3494_161 )
);
defparam \top/processor/sha_core/n3494_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [25]),
	.I2(\top/processor/sha_core/w[49] [25]),
	.F(\top/processor/sha_core/n3494_162 )
);
defparam \top/processor/sha_core/n3494_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [25]),
	.I2(\top/processor/sha_core/w[53] [25]),
	.F(\top/processor/sha_core/n3494_163 )
);
defparam \top/processor/sha_core/n3494_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_177 ),
	.I3(\top/processor/sha_core/n3494_162 ),
	.F(\top/processor/sha_core/n3866_124 )
);
defparam \top/processor/sha_core/n3866_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [25]),
	.I2(\top/processor/sha_core/w[55] [25]),
	.F(\top/processor/sha_core/n3866_125 )
);
defparam \top/processor/sha_core/n3866_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3618_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [20]),
	.I3(\top/processor/sha_core/w[37] [20]),
	.F(\top/processor/sha_core/n3618_165 )
);
defparam \top/processor/sha_core/n3618_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [19]),
	.I3(\top/processor/sha_core/w[37] [19]),
	.F(\top/processor/sha_core/n3619_165 )
);
defparam \top/processor/sha_core/n3619_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [18]),
	.I3(\top/processor/sha_core/w[37] [18]),
	.F(\top/processor/sha_core/n3620_165 )
);
defparam \top/processor/sha_core/n3620_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [17]),
	.I3(\top/processor/sha_core/w[37] [17]),
	.F(\top/processor/sha_core/n3621_165 )
);
defparam \top/processor/sha_core/n3621_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [16]),
	.I3(\top/processor/sha_core/w[37] [16]),
	.F(\top/processor/sha_core/n3622_165 )
);
defparam \top/processor/sha_core/n3622_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [15]),
	.I3(\top/processor/sha_core/w[37] [15]),
	.F(\top/processor/sha_core/n3623_165 )
);
defparam \top/processor/sha_core/n3623_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [14]),
	.I3(\top/processor/sha_core/w[37] [14]),
	.F(\top/processor/sha_core/n3624_165 )
);
defparam \top/processor/sha_core/n3624_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [13]),
	.I3(\top/processor/sha_core/w[37] [13]),
	.F(\top/processor/sha_core/n3625_165 )
);
defparam \top/processor/sha_core/n3625_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [12]),
	.I3(\top/processor/sha_core/w[37] [12]),
	.F(\top/processor/sha_core/n3626_165 )
);
defparam \top/processor/sha_core/n3626_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [11]),
	.I3(\top/processor/sha_core/w[37] [11]),
	.F(\top/processor/sha_core/n3627_165 )
);
defparam \top/processor/sha_core/n3627_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [10]),
	.I3(\top/processor/sha_core/w[37] [10]),
	.F(\top/processor/sha_core/n3628_165 )
);
defparam \top/processor/sha_core/n3628_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [9]),
	.I3(\top/processor/sha_core/w[37] [9]),
	.F(\top/processor/sha_core/n3629_165 )
);
defparam \top/processor/sha_core/n3629_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [8]),
	.I3(\top/processor/sha_core/w[37] [8]),
	.F(\top/processor/sha_core/n3630_165 )
);
defparam \top/processor/sha_core/n3630_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [7]),
	.I3(\top/processor/sha_core/w[37] [7]),
	.F(\top/processor/sha_core/n3631_165 )
);
defparam \top/processor/sha_core/n3631_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [6]),
	.I3(\top/processor/sha_core/w[37] [6]),
	.F(\top/processor/sha_core/n3632_165 )
);
defparam \top/processor/sha_core/n3632_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [5]),
	.I3(\top/processor/sha_core/w[37] [5]),
	.F(\top/processor/sha_core/n3633_165 )
);
defparam \top/processor/sha_core/n3633_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [4]),
	.I3(\top/processor/sha_core/w[37] [4]),
	.F(\top/processor/sha_core/n3634_165 )
);
defparam \top/processor/sha_core/n3634_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [3]),
	.I3(\top/processor/sha_core/w[37] [3]),
	.F(\top/processor/sha_core/n3635_165 )
);
defparam \top/processor/sha_core/n3635_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [2]),
	.I3(\top/processor/sha_core/w[37] [2]),
	.F(\top/processor/sha_core/n3636_165 )
);
defparam \top/processor/sha_core/n3636_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [1]),
	.I3(\top/processor/sha_core/w[37] [1]),
	.F(\top/processor/sha_core/n3637_165 )
);
defparam \top/processor/sha_core/n3637_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3494_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_127 ),
	.I3(\top/processor/sha_core/n3494_178 ),
	.F(\top/processor/sha_core/n3494_164 )
);
defparam \top/processor/sha_core/n3494_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [25]),
	.I2(\top/processor/sha_core/w[57] [25]),
	.F(\top/processor/sha_core/n3494_165 )
);
defparam \top/processor/sha_core/n3494_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [25]),
	.I2(\top/processor/sha_core/w[61] [25]),
	.F(\top/processor/sha_core/n3494_166 )
);
defparam \top/processor/sha_core/n3494_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_178 ),
	.I3(\top/processor/sha_core/n3494_165 ),
	.F(\top/processor/sha_core/n3866_126 )
);
defparam \top/processor/sha_core/n3866_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [25]),
	.I2(\top/processor/sha_core/w[63] [25]),
	.F(\top/processor/sha_core/n3866_127 )
);
defparam \top/processor/sha_core/n3866_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3638_s144  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[39] [0]),
	.I3(\top/processor/sha_core/w[37] [0]),
	.F(\top/processor/sha_core/n3638_165 )
);
defparam \top/processor/sha_core/n3638_s144 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_117 ),
	.I3(\top/processor/sha_core/n3495_172 ),
	.F(\top/processor/sha_core/n3495_148 )
);
defparam \top/processor/sha_core/n3495_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [24]),
	.I2(\top/processor/sha_core/w[1] [24]),
	.F(\top/processor/sha_core/n3495_149 )
);
defparam \top/processor/sha_core/n3495_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [24]),
	.I2(\top/processor/sha_core/w[5] [24]),
	.F(\top/processor/sha_core/n3495_150 )
);
defparam \top/processor/sha_core/n3495_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_172 ),
	.I3(\top/processor/sha_core/n3495_149 ),
	.F(\top/processor/sha_core/n3867_116 )
);
defparam \top/processor/sha_core/n3867_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [24]),
	.I2(\top/processor/sha_core/w[7] [24]),
	.F(\top/processor/sha_core/n3867_117 )
);
defparam \top/processor/sha_core/n3867_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [31]),
	.I3(\top/processor/sha_core/w[41] [31]),
	.F(\top/processor/sha_core/n3607_166 )
);
defparam \top/processor/sha_core/n3607_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [30]),
	.I3(\top/processor/sha_core/w[41] [30]),
	.F(\top/processor/sha_core/n3608_166 )
);
defparam \top/processor/sha_core/n3608_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [29]),
	.I3(\top/processor/sha_core/w[41] [29]),
	.F(\top/processor/sha_core/n3609_166 )
);
defparam \top/processor/sha_core/n3609_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [28]),
	.I3(\top/processor/sha_core/w[41] [28]),
	.F(\top/processor/sha_core/n3610_166 )
);
defparam \top/processor/sha_core/n3610_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [27]),
	.I3(\top/processor/sha_core/w[41] [27]),
	.F(\top/processor/sha_core/n3611_166 )
);
defparam \top/processor/sha_core/n3611_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [26]),
	.I3(\top/processor/sha_core/w[41] [26]),
	.F(\top/processor/sha_core/n3612_166 )
);
defparam \top/processor/sha_core/n3612_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [25]),
	.I3(\top/processor/sha_core/w[41] [25]),
	.F(\top/processor/sha_core/n3613_166 )
);
defparam \top/processor/sha_core/n3613_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_119 ),
	.I3(\top/processor/sha_core/n3495_173 ),
	.F(\top/processor/sha_core/n3495_151 )
);
defparam \top/processor/sha_core/n3495_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [24]),
	.I2(\top/processor/sha_core/w[9] [24]),
	.F(\top/processor/sha_core/n3495_152 )
);
defparam \top/processor/sha_core/n3495_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [24]),
	.I2(\top/processor/sha_core/w[13] [24]),
	.F(\top/processor/sha_core/n3495_153 )
);
defparam \top/processor/sha_core/n3495_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_173 ),
	.I3(\top/processor/sha_core/n3495_152 ),
	.F(\top/processor/sha_core/n3867_118 )
);
defparam \top/processor/sha_core/n3867_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [24]),
	.I2(\top/processor/sha_core/w[15] [24]),
	.F(\top/processor/sha_core/n3867_119 )
);
defparam \top/processor/sha_core/n3867_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3614_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [24]),
	.I3(\top/processor/sha_core/w[41] [24]),
	.F(\top/processor/sha_core/n3614_166 )
);
defparam \top/processor/sha_core/n3614_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [23]),
	.I3(\top/processor/sha_core/w[41] [23]),
	.F(\top/processor/sha_core/n3615_166 )
);
defparam \top/processor/sha_core/n3615_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [22]),
	.I3(\top/processor/sha_core/w[41] [22]),
	.F(\top/processor/sha_core/n3616_166 )
);
defparam \top/processor/sha_core/n3616_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [21]),
	.I3(\top/processor/sha_core/w[41] [21]),
	.F(\top/processor/sha_core/n3617_166 )
);
defparam \top/processor/sha_core/n3617_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [20]),
	.I3(\top/processor/sha_core/w[41] [20]),
	.F(\top/processor/sha_core/n3618_166 )
);
defparam \top/processor/sha_core/n3618_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [19]),
	.I3(\top/processor/sha_core/w[41] [19]),
	.F(\top/processor/sha_core/n3619_166 )
);
defparam \top/processor/sha_core/n3619_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [18]),
	.I3(\top/processor/sha_core/w[41] [18]),
	.F(\top/processor/sha_core/n3620_166 )
);
defparam \top/processor/sha_core/n3620_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [17]),
	.I3(\top/processor/sha_core/w[41] [17]),
	.F(\top/processor/sha_core/n3621_166 )
);
defparam \top/processor/sha_core/n3621_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [16]),
	.I3(\top/processor/sha_core/w[41] [16]),
	.F(\top/processor/sha_core/n3622_166 )
);
defparam \top/processor/sha_core/n3622_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [15]),
	.I3(\top/processor/sha_core/w[41] [15]),
	.F(\top/processor/sha_core/n3623_166 )
);
defparam \top/processor/sha_core/n3623_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [14]),
	.I3(\top/processor/sha_core/w[41] [14]),
	.F(\top/processor/sha_core/n3624_166 )
);
defparam \top/processor/sha_core/n3624_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [13]),
	.I3(\top/processor/sha_core/w[41] [13]),
	.F(\top/processor/sha_core/n3625_166 )
);
defparam \top/processor/sha_core/n3625_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [12]),
	.I3(\top/processor/sha_core/w[41] [12]),
	.F(\top/processor/sha_core/n3626_166 )
);
defparam \top/processor/sha_core/n3626_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [11]),
	.I3(\top/processor/sha_core/w[41] [11]),
	.F(\top/processor/sha_core/n3627_166 )
);
defparam \top/processor/sha_core/n3627_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [10]),
	.I3(\top/processor/sha_core/w[41] [10]),
	.F(\top/processor/sha_core/n3628_166 )
);
defparam \top/processor/sha_core/n3628_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [9]),
	.I3(\top/processor/sha_core/w[41] [9]),
	.F(\top/processor/sha_core/n3629_166 )
);
defparam \top/processor/sha_core/n3629_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [8]),
	.I3(\top/processor/sha_core/w[41] [8]),
	.F(\top/processor/sha_core/n3630_166 )
);
defparam \top/processor/sha_core/n3630_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [7]),
	.I3(\top/processor/sha_core/w[41] [7]),
	.F(\top/processor/sha_core/n3631_166 )
);
defparam \top/processor/sha_core/n3631_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [6]),
	.I3(\top/processor/sha_core/w[41] [6]),
	.F(\top/processor/sha_core/n3632_166 )
);
defparam \top/processor/sha_core/n3632_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [5]),
	.I3(\top/processor/sha_core/w[41] [5]),
	.F(\top/processor/sha_core/n3633_166 )
);
defparam \top/processor/sha_core/n3633_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_121 ),
	.I3(\top/processor/sha_core/n3495_174 ),
	.F(\top/processor/sha_core/n3495_154 )
);
defparam \top/processor/sha_core/n3495_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [24]),
	.I2(\top/processor/sha_core/w[17] [24]),
	.F(\top/processor/sha_core/n3495_155 )
);
defparam \top/processor/sha_core/n3495_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [24]),
	.I2(\top/processor/sha_core/w[21] [24]),
	.F(\top/processor/sha_core/n3495_156 )
);
defparam \top/processor/sha_core/n3495_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_174 ),
	.I3(\top/processor/sha_core/n3495_155 ),
	.F(\top/processor/sha_core/n3867_120 )
);
defparam \top/processor/sha_core/n3867_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [24]),
	.I2(\top/processor/sha_core/w[23] [24]),
	.F(\top/processor/sha_core/n3867_121 )
);
defparam \top/processor/sha_core/n3867_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3634_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [4]),
	.I3(\top/processor/sha_core/w[41] [4]),
	.F(\top/processor/sha_core/n3634_166 )
);
defparam \top/processor/sha_core/n3634_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [3]),
	.I3(\top/processor/sha_core/w[41] [3]),
	.F(\top/processor/sha_core/n3635_166 )
);
defparam \top/processor/sha_core/n3635_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [2]),
	.I3(\top/processor/sha_core/w[41] [2]),
	.F(\top/processor/sha_core/n3636_166 )
);
defparam \top/processor/sha_core/n3636_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [1]),
	.I3(\top/processor/sha_core/w[41] [1]),
	.F(\top/processor/sha_core/n3637_166 )
);
defparam \top/processor/sha_core/n3637_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[43] [0]),
	.I3(\top/processor/sha_core/w[41] [0]),
	.F(\top/processor/sha_core/n3638_166 )
);
defparam \top/processor/sha_core/n3638_s145 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_123 ),
	.I3(\top/processor/sha_core/n3495_175 ),
	.F(\top/processor/sha_core/n3495_157 )
);
defparam \top/processor/sha_core/n3495_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [24]),
	.I2(\top/processor/sha_core/w[25] [24]),
	.F(\top/processor/sha_core/n3495_158 )
);
defparam \top/processor/sha_core/n3495_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [24]),
	.I2(\top/processor/sha_core/w[29] [24]),
	.F(\top/processor/sha_core/n3495_159 )
);
defparam \top/processor/sha_core/n3495_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_175 ),
	.I3(\top/processor/sha_core/n3495_158 ),
	.F(\top/processor/sha_core/n3867_122 )
);
defparam \top/processor/sha_core/n3867_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [24]),
	.I2(\top/processor/sha_core/w[31] [24]),
	.F(\top/processor/sha_core/n3867_123 )
);
defparam \top/processor/sha_core/n3867_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_117 ),
	.I3(\top/processor/sha_core/n3488_172 ),
	.F(\top/processor/sha_core/n3488_148 )
);
defparam \top/processor/sha_core/n3488_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [31]),
	.I2(\top/processor/sha_core/w[41] [31]),
	.F(\top/processor/sha_core/n3488_149 )
);
defparam \top/processor/sha_core/n3488_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [31]),
	.I2(\top/processor/sha_core/w[45] [31]),
	.F(\top/processor/sha_core/n3488_150 )
);
defparam \top/processor/sha_core/n3488_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_172 ),
	.I3(\top/processor/sha_core/n3488_149 ),
	.F(\top/processor/sha_core/n3860_116 )
);
defparam \top/processor/sha_core/n3860_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [31]),
	.I2(\top/processor/sha_core/w[47] [31]),
	.F(\top/processor/sha_core/n3860_117 )
);
defparam \top/processor/sha_core/n3860_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [31]),
	.I3(\top/processor/sha_core/w[45] [31]),
	.F(\top/processor/sha_core/n3607_167 )
);
defparam \top/processor/sha_core/n3607_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [30]),
	.I3(\top/processor/sha_core/w[45] [30]),
	.F(\top/processor/sha_core/n3608_167 )
);
defparam \top/processor/sha_core/n3608_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [29]),
	.I3(\top/processor/sha_core/w[45] [29]),
	.F(\top/processor/sha_core/n3609_167 )
);
defparam \top/processor/sha_core/n3609_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_125 ),
	.I3(\top/processor/sha_core/n3495_176 ),
	.F(\top/processor/sha_core/n3495_160 )
);
defparam \top/processor/sha_core/n3495_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [24]),
	.I2(\top/processor/sha_core/w[33] [24]),
	.F(\top/processor/sha_core/n3495_161 )
);
defparam \top/processor/sha_core/n3495_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [24]),
	.I2(\top/processor/sha_core/w[37] [24]),
	.F(\top/processor/sha_core/n3495_162 )
);
defparam \top/processor/sha_core/n3495_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_176 ),
	.I3(\top/processor/sha_core/n3495_161 ),
	.F(\top/processor/sha_core/n3867_124 )
);
defparam \top/processor/sha_core/n3867_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [24]),
	.I2(\top/processor/sha_core/w[39] [24]),
	.F(\top/processor/sha_core/n3867_125 )
);
defparam \top/processor/sha_core/n3867_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3610_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [28]),
	.I3(\top/processor/sha_core/w[45] [28]),
	.F(\top/processor/sha_core/n3610_167 )
);
defparam \top/processor/sha_core/n3610_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [27]),
	.I3(\top/processor/sha_core/w[45] [27]),
	.F(\top/processor/sha_core/n3611_167 )
);
defparam \top/processor/sha_core/n3611_s146 .INIT=16'hD9C8;
LUT4 \top/processor/sha_core/n3612_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [26]),
	.I3(\top/processor/sha_core/w[45] [26]),
	.F(\top/processor/sha_core/n3612_167 )
);
defparam \top/processor/sha_core/n3612_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [25]),
	.I3(\top/processor/sha_core/w[45] [25]),
	.F(\top/processor/sha_core/n3613_167 )
);
defparam \top/processor/sha_core/n3613_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [24]),
	.I3(\top/processor/sha_core/w[45] [24]),
	.F(\top/processor/sha_core/n3614_167 )
);
defparam \top/processor/sha_core/n3614_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [23]),
	.I3(\top/processor/sha_core/w[45] [23]),
	.F(\top/processor/sha_core/n3615_167 )
);
defparam \top/processor/sha_core/n3615_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [22]),
	.I3(\top/processor/sha_core/w[45] [22]),
	.F(\top/processor/sha_core/n3616_167 )
);
defparam \top/processor/sha_core/n3616_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [21]),
	.I3(\top/processor/sha_core/w[45] [21]),
	.F(\top/processor/sha_core/n3617_167 )
);
defparam \top/processor/sha_core/n3617_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [20]),
	.I3(\top/processor/sha_core/w[45] [20]),
	.F(\top/processor/sha_core/n3618_167 )
);
defparam \top/processor/sha_core/n3618_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [19]),
	.I3(\top/processor/sha_core/w[45] [19]),
	.F(\top/processor/sha_core/n3619_167 )
);
defparam \top/processor/sha_core/n3619_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [18]),
	.I3(\top/processor/sha_core/w[45] [18]),
	.F(\top/processor/sha_core/n3620_167 )
);
defparam \top/processor/sha_core/n3620_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [17]),
	.I3(\top/processor/sha_core/w[45] [17]),
	.F(\top/processor/sha_core/n3621_167 )
);
defparam \top/processor/sha_core/n3621_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [16]),
	.I3(\top/processor/sha_core/w[45] [16]),
	.F(\top/processor/sha_core/n3622_167 )
);
defparam \top/processor/sha_core/n3622_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [15]),
	.I3(\top/processor/sha_core/w[45] [15]),
	.F(\top/processor/sha_core/n3623_167 )
);
defparam \top/processor/sha_core/n3623_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [14]),
	.I3(\top/processor/sha_core/w[45] [14]),
	.F(\top/processor/sha_core/n3624_167 )
);
defparam \top/processor/sha_core/n3624_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [13]),
	.I3(\top/processor/sha_core/w[45] [13]),
	.F(\top/processor/sha_core/n3625_167 )
);
defparam \top/processor/sha_core/n3625_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [12]),
	.I3(\top/processor/sha_core/w[45] [12]),
	.F(\top/processor/sha_core/n3626_167 )
);
defparam \top/processor/sha_core/n3626_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [11]),
	.I3(\top/processor/sha_core/w[45] [11]),
	.F(\top/processor/sha_core/n3627_167 )
);
defparam \top/processor/sha_core/n3627_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [10]),
	.I3(\top/processor/sha_core/w[45] [10]),
	.F(\top/processor/sha_core/n3628_167 )
);
defparam \top/processor/sha_core/n3628_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [9]),
	.I3(\top/processor/sha_core/w[45] [9]),
	.F(\top/processor/sha_core/n3629_167 )
);
defparam \top/processor/sha_core/n3629_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_127 ),
	.I3(\top/processor/sha_core/n3495_177 ),
	.F(\top/processor/sha_core/n3495_163 )
);
defparam \top/processor/sha_core/n3495_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [24]),
	.I2(\top/processor/sha_core/w[41] [24]),
	.F(\top/processor/sha_core/n3495_164 )
);
defparam \top/processor/sha_core/n3495_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [24]),
	.I2(\top/processor/sha_core/w[45] [24]),
	.F(\top/processor/sha_core/n3495_165 )
);
defparam \top/processor/sha_core/n3495_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_177 ),
	.I3(\top/processor/sha_core/n3495_164 ),
	.F(\top/processor/sha_core/n3867_126 )
);
defparam \top/processor/sha_core/n3867_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [24]),
	.I2(\top/processor/sha_core/w[47] [24]),
	.F(\top/processor/sha_core/n3867_127 )
);
defparam \top/processor/sha_core/n3867_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3630_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [8]),
	.I3(\top/processor/sha_core/w[45] [8]),
	.F(\top/processor/sha_core/n3630_167 )
);
defparam \top/processor/sha_core/n3630_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [7]),
	.I3(\top/processor/sha_core/w[45] [7]),
	.F(\top/processor/sha_core/n3631_167 )
);
defparam \top/processor/sha_core/n3631_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [6]),
	.I3(\top/processor/sha_core/w[45] [6]),
	.F(\top/processor/sha_core/n3632_167 )
);
defparam \top/processor/sha_core/n3632_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [5]),
	.I3(\top/processor/sha_core/w[45] [5]),
	.F(\top/processor/sha_core/n3633_167 )
);
defparam \top/processor/sha_core/n3633_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [4]),
	.I3(\top/processor/sha_core/w[45] [4]),
	.F(\top/processor/sha_core/n3634_167 )
);
defparam \top/processor/sha_core/n3634_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [3]),
	.I3(\top/processor/sha_core/w[45] [3]),
	.F(\top/processor/sha_core/n3635_167 )
);
defparam \top/processor/sha_core/n3635_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [2]),
	.I3(\top/processor/sha_core/w[45] [2]),
	.F(\top/processor/sha_core/n3636_167 )
);
defparam \top/processor/sha_core/n3636_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [1]),
	.I3(\top/processor/sha_core/w[45] [1]),
	.F(\top/processor/sha_core/n3637_167 )
);
defparam \top/processor/sha_core/n3637_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[47] [0]),
	.I3(\top/processor/sha_core/w[45] [0]),
	.F(\top/processor/sha_core/n3638_167 )
);
defparam \top/processor/sha_core/n3638_s146 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3495_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_129 ),
	.I3(\top/processor/sha_core/n3495_178 ),
	.F(\top/processor/sha_core/n3495_166 )
);
defparam \top/processor/sha_core/n3495_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [24]),
	.I2(\top/processor/sha_core/w[49] [24]),
	.F(\top/processor/sha_core/n3495_167 )
);
defparam \top/processor/sha_core/n3495_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [24]),
	.I2(\top/processor/sha_core/w[53] [24]),
	.F(\top/processor/sha_core/n3495_168 )
);
defparam \top/processor/sha_core/n3495_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_178 ),
	.I3(\top/processor/sha_core/n3495_167 ),
	.F(\top/processor/sha_core/n3867_128 )
);
defparam \top/processor/sha_core/n3867_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [24]),
	.I2(\top/processor/sha_core/w[55] [24]),
	.F(\top/processor/sha_core/n3867_129 )
);
defparam \top/processor/sha_core/n3867_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3495_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3867_131 ),
	.I3(\top/processor/sha_core/n3495_179 ),
	.F(\top/processor/sha_core/n3495_169 )
);
defparam \top/processor/sha_core/n3495_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3495_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [24]),
	.I2(\top/processor/sha_core/w[57] [24]),
	.F(\top/processor/sha_core/n3495_170 )
);
defparam \top/processor/sha_core/n3495_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [24]),
	.I2(\top/processor/sha_core/w[61] [24]),
	.F(\top/processor/sha_core/n3495_171 )
);
defparam \top/processor/sha_core/n3495_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3867_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3495_179 ),
	.I3(\top/processor/sha_core/n3495_170 ),
	.F(\top/processor/sha_core/n3867_130 )
);
defparam \top/processor/sha_core/n3867_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3867_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [24]),
	.I2(\top/processor/sha_core/w[63] [24]),
	.F(\top/processor/sha_core/n3867_131 )
);
defparam \top/processor/sha_core/n3867_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [31]),
	.I3(\top/processor/sha_core/w[49] [31]),
	.F(\top/processor/sha_core/n3607_168 )
);
defparam \top/processor/sha_core/n3607_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [30]),
	.I3(\top/processor/sha_core/w[49] [30]),
	.F(\top/processor/sha_core/n3608_168 )
);
defparam \top/processor/sha_core/n3608_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [29]),
	.I3(\top/processor/sha_core/w[49] [29]),
	.F(\top/processor/sha_core/n3609_168 )
);
defparam \top/processor/sha_core/n3609_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [28]),
	.I3(\top/processor/sha_core/w[49] [28]),
	.F(\top/processor/sha_core/n3610_168 )
);
defparam \top/processor/sha_core/n3610_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [27]),
	.I3(\top/processor/sha_core/w[49] [27]),
	.F(\top/processor/sha_core/n3611_168 )
);
defparam \top/processor/sha_core/n3611_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [26]),
	.I3(\top/processor/sha_core/w[49] [26]),
	.F(\top/processor/sha_core/n3612_168 )
);
defparam \top/processor/sha_core/n3612_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [25]),
	.I3(\top/processor/sha_core/w[49] [25]),
	.F(\top/processor/sha_core/n3613_168 )
);
defparam \top/processor/sha_core/n3613_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [24]),
	.I3(\top/processor/sha_core/w[49] [24]),
	.F(\top/processor/sha_core/n3614_168 )
);
defparam \top/processor/sha_core/n3614_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [23]),
	.I3(\top/processor/sha_core/w[49] [23]),
	.F(\top/processor/sha_core/n3615_168 )
);
defparam \top/processor/sha_core/n3615_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [22]),
	.I3(\top/processor/sha_core/w[49] [22]),
	.F(\top/processor/sha_core/n3616_168 )
);
defparam \top/processor/sha_core/n3616_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [21]),
	.I3(\top/processor/sha_core/w[49] [21]),
	.F(\top/processor/sha_core/n3617_168 )
);
defparam \top/processor/sha_core/n3617_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [20]),
	.I3(\top/processor/sha_core/w[49] [20]),
	.F(\top/processor/sha_core/n3618_168 )
);
defparam \top/processor/sha_core/n3618_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [19]),
	.I3(\top/processor/sha_core/w[49] [19]),
	.F(\top/processor/sha_core/n3619_168 )
);
defparam \top/processor/sha_core/n3619_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [18]),
	.I3(\top/processor/sha_core/w[49] [18]),
	.F(\top/processor/sha_core/n3620_168 )
);
defparam \top/processor/sha_core/n3620_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [17]),
	.I3(\top/processor/sha_core/w[49] [17]),
	.F(\top/processor/sha_core/n3621_168 )
);
defparam \top/processor/sha_core/n3621_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [16]),
	.I3(\top/processor/sha_core/w[49] [16]),
	.F(\top/processor/sha_core/n3622_168 )
);
defparam \top/processor/sha_core/n3622_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [15]),
	.I3(\top/processor/sha_core/w[49] [15]),
	.F(\top/processor/sha_core/n3623_168 )
);
defparam \top/processor/sha_core/n3623_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [14]),
	.I3(\top/processor/sha_core/w[49] [14]),
	.F(\top/processor/sha_core/n3624_168 )
);
defparam \top/processor/sha_core/n3624_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [13]),
	.I3(\top/processor/sha_core/w[49] [13]),
	.F(\top/processor/sha_core/n3625_168 )
);
defparam \top/processor/sha_core/n3625_s147 .INIT=16'hD9C8;
LUT4 \top/processor/sha_core/n3496_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_117 ),
	.I3(\top/processor/sha_core/n3496_172 ),
	.F(\top/processor/sha_core/n3496_148 )
);
defparam \top/processor/sha_core/n3496_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [23]),
	.I2(\top/processor/sha_core/w[1] [23]),
	.F(\top/processor/sha_core/n3496_149 )
);
defparam \top/processor/sha_core/n3496_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [23]),
	.I2(\top/processor/sha_core/w[5] [23]),
	.F(\top/processor/sha_core/n3496_150 )
);
defparam \top/processor/sha_core/n3496_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_172 ),
	.I3(\top/processor/sha_core/n3496_149 ),
	.F(\top/processor/sha_core/n3868_116 )
);
defparam \top/processor/sha_core/n3868_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [23]),
	.I2(\top/processor/sha_core/w[7] [23]),
	.F(\top/processor/sha_core/n3868_117 )
);
defparam \top/processor/sha_core/n3868_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3626_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [12]),
	.I3(\top/processor/sha_core/w[49] [12]),
	.F(\top/processor/sha_core/n3626_168 )
);
defparam \top/processor/sha_core/n3626_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [11]),
	.I3(\top/processor/sha_core/w[49] [11]),
	.F(\top/processor/sha_core/n3627_168 )
);
defparam \top/processor/sha_core/n3627_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [10]),
	.I3(\top/processor/sha_core/w[49] [10]),
	.F(\top/processor/sha_core/n3628_168 )
);
defparam \top/processor/sha_core/n3628_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [9]),
	.I3(\top/processor/sha_core/w[49] [9]),
	.F(\top/processor/sha_core/n3629_168 )
);
defparam \top/processor/sha_core/n3629_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [8]),
	.I3(\top/processor/sha_core/w[49] [8]),
	.F(\top/processor/sha_core/n3630_168 )
);
defparam \top/processor/sha_core/n3630_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [7]),
	.I3(\top/processor/sha_core/w[49] [7]),
	.F(\top/processor/sha_core/n3631_168 )
);
defparam \top/processor/sha_core/n3631_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [6]),
	.I3(\top/processor/sha_core/w[49] [6]),
	.F(\top/processor/sha_core/n3632_168 )
);
defparam \top/processor/sha_core/n3632_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [5]),
	.I3(\top/processor/sha_core/w[49] [5]),
	.F(\top/processor/sha_core/n3633_168 )
);
defparam \top/processor/sha_core/n3633_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [4]),
	.I3(\top/processor/sha_core/w[49] [4]),
	.F(\top/processor/sha_core/n3634_168 )
);
defparam \top/processor/sha_core/n3634_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [3]),
	.I3(\top/processor/sha_core/w[49] [3]),
	.F(\top/processor/sha_core/n3635_168 )
);
defparam \top/processor/sha_core/n3635_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [2]),
	.I3(\top/processor/sha_core/w[49] [2]),
	.F(\top/processor/sha_core/n3636_168 )
);
defparam \top/processor/sha_core/n3636_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [1]),
	.I3(\top/processor/sha_core/w[49] [1]),
	.F(\top/processor/sha_core/n3637_168 )
);
defparam \top/processor/sha_core/n3637_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s147  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[51] [0]),
	.I3(\top/processor/sha_core/w[49] [0]),
	.F(\top/processor/sha_core/n3638_168 )
);
defparam \top/processor/sha_core/n3638_s147 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3496_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_119 ),
	.I3(\top/processor/sha_core/n3496_173 ),
	.F(\top/processor/sha_core/n3496_151 )
);
defparam \top/processor/sha_core/n3496_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [23]),
	.I2(\top/processor/sha_core/w[9] [23]),
	.F(\top/processor/sha_core/n3496_152 )
);
defparam \top/processor/sha_core/n3496_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [23]),
	.I2(\top/processor/sha_core/w[13] [23]),
	.F(\top/processor/sha_core/n3496_153 )
);
defparam \top/processor/sha_core/n3496_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_173 ),
	.I3(\top/processor/sha_core/n3496_152 ),
	.F(\top/processor/sha_core/n3868_118 )
);
defparam \top/processor/sha_core/n3868_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [23]),
	.I2(\top/processor/sha_core/w[15] [23]),
	.F(\top/processor/sha_core/n3868_119 )
);
defparam \top/processor/sha_core/n3868_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3496_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_121 ),
	.I3(\top/processor/sha_core/n3496_174 ),
	.F(\top/processor/sha_core/n3496_154 )
);
defparam \top/processor/sha_core/n3496_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [23]),
	.I2(\top/processor/sha_core/w[17] [23]),
	.F(\top/processor/sha_core/n3496_155 )
);
defparam \top/processor/sha_core/n3496_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [23]),
	.I2(\top/processor/sha_core/w[21] [23]),
	.F(\top/processor/sha_core/n3496_156 )
);
defparam \top/processor/sha_core/n3496_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_174 ),
	.I3(\top/processor/sha_core/n3496_155 ),
	.F(\top/processor/sha_core/n3868_120 )
);
defparam \top/processor/sha_core/n3868_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [23]),
	.I2(\top/processor/sha_core/w[23] [23]),
	.F(\top/processor/sha_core/n3868_121 )
);
defparam \top/processor/sha_core/n3868_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [31]),
	.I3(\top/processor/sha_core/w[53] [31]),
	.F(\top/processor/sha_core/n3607_169 )
);
defparam \top/processor/sha_core/n3607_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [30]),
	.I3(\top/processor/sha_core/w[53] [30]),
	.F(\top/processor/sha_core/n3608_169 )
);
defparam \top/processor/sha_core/n3608_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [29]),
	.I3(\top/processor/sha_core/w[53] [29]),
	.F(\top/processor/sha_core/n3609_169 )
);
defparam \top/processor/sha_core/n3609_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [28]),
	.I3(\top/processor/sha_core/w[53] [28]),
	.F(\top/processor/sha_core/n3610_169 )
);
defparam \top/processor/sha_core/n3610_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [27]),
	.I3(\top/processor/sha_core/w[53] [27]),
	.F(\top/processor/sha_core/n3611_169 )
);
defparam \top/processor/sha_core/n3611_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [26]),
	.I3(\top/processor/sha_core/w[53] [26]),
	.F(\top/processor/sha_core/n3612_169 )
);
defparam \top/processor/sha_core/n3612_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [25]),
	.I3(\top/processor/sha_core/w[53] [25]),
	.F(\top/processor/sha_core/n3613_169 )
);
defparam \top/processor/sha_core/n3613_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [24]),
	.I3(\top/processor/sha_core/w[53] [24]),
	.F(\top/processor/sha_core/n3614_169 )
);
defparam \top/processor/sha_core/n3614_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [23]),
	.I3(\top/processor/sha_core/w[53] [23]),
	.F(\top/processor/sha_core/n3615_169 )
);
defparam \top/processor/sha_core/n3615_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [22]),
	.I3(\top/processor/sha_core/w[53] [22]),
	.F(\top/processor/sha_core/n3616_169 )
);
defparam \top/processor/sha_core/n3616_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [21]),
	.I3(\top/processor/sha_core/w[53] [21]),
	.F(\top/processor/sha_core/n3617_169 )
);
defparam \top/processor/sha_core/n3617_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [20]),
	.I3(\top/processor/sha_core/w[53] [20]),
	.F(\top/processor/sha_core/n3618_169 )
);
defparam \top/processor/sha_core/n3618_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [19]),
	.I3(\top/processor/sha_core/w[53] [19]),
	.F(\top/processor/sha_core/n3619_169 )
);
defparam \top/processor/sha_core/n3619_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [18]),
	.I3(\top/processor/sha_core/w[53] [18]),
	.F(\top/processor/sha_core/n3620_169 )
);
defparam \top/processor/sha_core/n3620_s148 .INIT=16'hD9C8;
LUT4 \top/processor/sha_core/n3621_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [17]),
	.I3(\top/processor/sha_core/w[53] [17]),
	.F(\top/processor/sha_core/n3621_169 )
);
defparam \top/processor/sha_core/n3621_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3496_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_123 ),
	.I3(\top/processor/sha_core/n3496_175 ),
	.F(\top/processor/sha_core/n3496_157 )
);
defparam \top/processor/sha_core/n3496_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [23]),
	.I2(\top/processor/sha_core/w[25] [23]),
	.F(\top/processor/sha_core/n3496_158 )
);
defparam \top/processor/sha_core/n3496_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [23]),
	.I2(\top/processor/sha_core/w[29] [23]),
	.F(\top/processor/sha_core/n3496_159 )
);
defparam \top/processor/sha_core/n3496_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_175 ),
	.I3(\top/processor/sha_core/n3496_158 ),
	.F(\top/processor/sha_core/n3868_122 )
);
defparam \top/processor/sha_core/n3868_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [23]),
	.I2(\top/processor/sha_core/w[31] [23]),
	.F(\top/processor/sha_core/n3868_123 )
);
defparam \top/processor/sha_core/n3868_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3622_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [16]),
	.I3(\top/processor/sha_core/w[53] [16]),
	.F(\top/processor/sha_core/n3622_169 )
);
defparam \top/processor/sha_core/n3622_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [15]),
	.I3(\top/processor/sha_core/w[53] [15]),
	.F(\top/processor/sha_core/n3623_169 )
);
defparam \top/processor/sha_core/n3623_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [14]),
	.I3(\top/processor/sha_core/w[53] [14]),
	.F(\top/processor/sha_core/n3624_169 )
);
defparam \top/processor/sha_core/n3624_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [13]),
	.I3(\top/processor/sha_core/w[53] [13]),
	.F(\top/processor/sha_core/n3625_169 )
);
defparam \top/processor/sha_core/n3625_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [12]),
	.I3(\top/processor/sha_core/w[53] [12]),
	.F(\top/processor/sha_core/n3626_169 )
);
defparam \top/processor/sha_core/n3626_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [11]),
	.I3(\top/processor/sha_core/w[53] [11]),
	.F(\top/processor/sha_core/n3627_169 )
);
defparam \top/processor/sha_core/n3627_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [10]),
	.I3(\top/processor/sha_core/w[53] [10]),
	.F(\top/processor/sha_core/n3628_169 )
);
defparam \top/processor/sha_core/n3628_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [9]),
	.I3(\top/processor/sha_core/w[53] [9]),
	.F(\top/processor/sha_core/n3629_169 )
);
defparam \top/processor/sha_core/n3629_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [8]),
	.I3(\top/processor/sha_core/w[53] [8]),
	.F(\top/processor/sha_core/n3630_169 )
);
defparam \top/processor/sha_core/n3630_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [7]),
	.I3(\top/processor/sha_core/w[53] [7]),
	.F(\top/processor/sha_core/n3631_169 )
);
defparam \top/processor/sha_core/n3631_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [6]),
	.I3(\top/processor/sha_core/w[53] [6]),
	.F(\top/processor/sha_core/n3632_169 )
);
defparam \top/processor/sha_core/n3632_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [5]),
	.I3(\top/processor/sha_core/w[53] [5]),
	.F(\top/processor/sha_core/n3633_169 )
);
defparam \top/processor/sha_core/n3633_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [4]),
	.I3(\top/processor/sha_core/w[53] [4]),
	.F(\top/processor/sha_core/n3634_169 )
);
defparam \top/processor/sha_core/n3634_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [3]),
	.I3(\top/processor/sha_core/w[53] [3]),
	.F(\top/processor/sha_core/n3635_169 )
);
defparam \top/processor/sha_core/n3635_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [2]),
	.I3(\top/processor/sha_core/w[53] [2]),
	.F(\top/processor/sha_core/n3636_169 )
);
defparam \top/processor/sha_core/n3636_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [1]),
	.I3(\top/processor/sha_core/w[53] [1]),
	.F(\top/processor/sha_core/n3637_169 )
);
defparam \top/processor/sha_core/n3637_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[55] [0]),
	.I3(\top/processor/sha_core/w[53] [0]),
	.F(\top/processor/sha_core/n3638_169 )
);
defparam \top/processor/sha_core/n3638_s148 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3496_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_125 ),
	.I3(\top/processor/sha_core/n3496_176 ),
	.F(\top/processor/sha_core/n3496_160 )
);
defparam \top/processor/sha_core/n3496_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [23]),
	.I2(\top/processor/sha_core/w[33] [23]),
	.F(\top/processor/sha_core/n3496_161 )
);
defparam \top/processor/sha_core/n3496_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [23]),
	.I2(\top/processor/sha_core/w[37] [23]),
	.F(\top/processor/sha_core/n3496_162 )
);
defparam \top/processor/sha_core/n3496_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_176 ),
	.I3(\top/processor/sha_core/n3496_161 ),
	.F(\top/processor/sha_core/n3868_124 )
);
defparam \top/processor/sha_core/n3868_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [23]),
	.I2(\top/processor/sha_core/w[39] [23]),
	.F(\top/processor/sha_core/n3868_125 )
);
defparam \top/processor/sha_core/n3868_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3496_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_127 ),
	.I3(\top/processor/sha_core/n3496_177 ),
	.F(\top/processor/sha_core/n3496_163 )
);
defparam \top/processor/sha_core/n3496_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [23]),
	.I2(\top/processor/sha_core/w[41] [23]),
	.F(\top/processor/sha_core/n3496_164 )
);
defparam \top/processor/sha_core/n3496_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [23]),
	.I2(\top/processor/sha_core/w[45] [23]),
	.F(\top/processor/sha_core/n3496_165 )
);
defparam \top/processor/sha_core/n3496_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_177 ),
	.I3(\top/processor/sha_core/n3496_164 ),
	.F(\top/processor/sha_core/n3868_126 )
);
defparam \top/processor/sha_core/n3868_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [23]),
	.I2(\top/processor/sha_core/w[47] [23]),
	.F(\top/processor/sha_core/n3868_127 )
);
defparam \top/processor/sha_core/n3868_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_119 ),
	.I3(\top/processor/sha_core/n3488_173 ),
	.F(\top/processor/sha_core/n3488_151 )
);
defparam \top/processor/sha_core/n3488_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [31]),
	.I2(\top/processor/sha_core/w[49] [31]),
	.F(\top/processor/sha_core/n3488_152 )
);
defparam \top/processor/sha_core/n3488_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [31]),
	.I2(\top/processor/sha_core/w[53] [31]),
	.F(\top/processor/sha_core/n3488_153 )
);
defparam \top/processor/sha_core/n3488_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_173 ),
	.I3(\top/processor/sha_core/n3488_152 ),
	.F(\top/processor/sha_core/n3860_118 )
);
defparam \top/processor/sha_core/n3860_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [31]),
	.I2(\top/processor/sha_core/w[55] [31]),
	.F(\top/processor/sha_core/n3860_119 )
);
defparam \top/processor/sha_core/n3860_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [31]),
	.I3(\top/processor/sha_core/w[57] [31]),
	.F(\top/processor/sha_core/n3607_170 )
);
defparam \top/processor/sha_core/n3607_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [30]),
	.I3(\top/processor/sha_core/w[57] [30]),
	.F(\top/processor/sha_core/n3608_170 )
);
defparam \top/processor/sha_core/n3608_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [29]),
	.I3(\top/processor/sha_core/w[57] [29]),
	.F(\top/processor/sha_core/n3609_170 )
);
defparam \top/processor/sha_core/n3609_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [28]),
	.I3(\top/processor/sha_core/w[57] [28]),
	.F(\top/processor/sha_core/n3610_170 )
);
defparam \top/processor/sha_core/n3610_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [27]),
	.I3(\top/processor/sha_core/w[57] [27]),
	.F(\top/processor/sha_core/n3611_170 )
);
defparam \top/processor/sha_core/n3611_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [26]),
	.I3(\top/processor/sha_core/w[57] [26]),
	.F(\top/processor/sha_core/n3612_170 )
);
defparam \top/processor/sha_core/n3612_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [25]),
	.I3(\top/processor/sha_core/w[57] [25]),
	.F(\top/processor/sha_core/n3613_170 )
);
defparam \top/processor/sha_core/n3613_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [24]),
	.I3(\top/processor/sha_core/w[57] [24]),
	.F(\top/processor/sha_core/n3614_170 )
);
defparam \top/processor/sha_core/n3614_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [23]),
	.I3(\top/processor/sha_core/w[57] [23]),
	.F(\top/processor/sha_core/n3615_170 )
);
defparam \top/processor/sha_core/n3615_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [22]),
	.I3(\top/processor/sha_core/w[57] [22]),
	.F(\top/processor/sha_core/n3616_170 )
);
defparam \top/processor/sha_core/n3616_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [21]),
	.I3(\top/processor/sha_core/w[57] [21]),
	.F(\top/processor/sha_core/n3617_170 )
);
defparam \top/processor/sha_core/n3617_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3496_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_129 ),
	.I3(\top/processor/sha_core/n3496_178 ),
	.F(\top/processor/sha_core/n3496_166 )
);
defparam \top/processor/sha_core/n3496_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [23]),
	.I2(\top/processor/sha_core/w[49] [23]),
	.F(\top/processor/sha_core/n3496_167 )
);
defparam \top/processor/sha_core/n3496_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [23]),
	.I2(\top/processor/sha_core/w[53] [23]),
	.F(\top/processor/sha_core/n3496_168 )
);
defparam \top/processor/sha_core/n3496_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_178 ),
	.I3(\top/processor/sha_core/n3496_167 ),
	.F(\top/processor/sha_core/n3868_128 )
);
defparam \top/processor/sha_core/n3868_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [23]),
	.I2(\top/processor/sha_core/w[55] [23]),
	.F(\top/processor/sha_core/n3868_129 )
);
defparam \top/processor/sha_core/n3868_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3618_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [20]),
	.I3(\top/processor/sha_core/w[57] [20]),
	.F(\top/processor/sha_core/n3618_170 )
);
defparam \top/processor/sha_core/n3618_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [19]),
	.I3(\top/processor/sha_core/w[57] [19]),
	.F(\top/processor/sha_core/n3619_170 )
);
defparam \top/processor/sha_core/n3619_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [18]),
	.I3(\top/processor/sha_core/w[57] [18]),
	.F(\top/processor/sha_core/n3620_170 )
);
defparam \top/processor/sha_core/n3620_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [17]),
	.I3(\top/processor/sha_core/w[57] [17]),
	.F(\top/processor/sha_core/n3621_170 )
);
defparam \top/processor/sha_core/n3621_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [16]),
	.I3(\top/processor/sha_core/w[57] [16]),
	.F(\top/processor/sha_core/n3622_170 )
);
defparam \top/processor/sha_core/n3622_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [15]),
	.I3(\top/processor/sha_core/w[57] [15]),
	.F(\top/processor/sha_core/n3623_170 )
);
defparam \top/processor/sha_core/n3623_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [14]),
	.I3(\top/processor/sha_core/w[57] [14]),
	.F(\top/processor/sha_core/n3624_170 )
);
defparam \top/processor/sha_core/n3624_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [13]),
	.I3(\top/processor/sha_core/w[57] [13]),
	.F(\top/processor/sha_core/n3625_170 )
);
defparam \top/processor/sha_core/n3625_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [12]),
	.I3(\top/processor/sha_core/w[57] [12]),
	.F(\top/processor/sha_core/n3626_170 )
);
defparam \top/processor/sha_core/n3626_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [11]),
	.I3(\top/processor/sha_core/w[57] [11]),
	.F(\top/processor/sha_core/n3627_170 )
);
defparam \top/processor/sha_core/n3627_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [10]),
	.I3(\top/processor/sha_core/w[57] [10]),
	.F(\top/processor/sha_core/n3628_170 )
);
defparam \top/processor/sha_core/n3628_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [9]),
	.I3(\top/processor/sha_core/w[57] [9]),
	.F(\top/processor/sha_core/n3629_170 )
);
defparam \top/processor/sha_core/n3629_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [8]),
	.I3(\top/processor/sha_core/w[57] [8]),
	.F(\top/processor/sha_core/n3630_170 )
);
defparam \top/processor/sha_core/n3630_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [7]),
	.I3(\top/processor/sha_core/w[57] [7]),
	.F(\top/processor/sha_core/n3631_170 )
);
defparam \top/processor/sha_core/n3631_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [6]),
	.I3(\top/processor/sha_core/w[57] [6]),
	.F(\top/processor/sha_core/n3632_170 )
);
defparam \top/processor/sha_core/n3632_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [5]),
	.I3(\top/processor/sha_core/w[57] [5]),
	.F(\top/processor/sha_core/n3633_170 )
);
defparam \top/processor/sha_core/n3633_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [4]),
	.I3(\top/processor/sha_core/w[57] [4]),
	.F(\top/processor/sha_core/n3634_170 )
);
defparam \top/processor/sha_core/n3634_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [3]),
	.I3(\top/processor/sha_core/w[57] [3]),
	.F(\top/processor/sha_core/n3635_170 )
);
defparam \top/processor/sha_core/n3635_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [2]),
	.I3(\top/processor/sha_core/w[57] [2]),
	.F(\top/processor/sha_core/n3636_170 )
);
defparam \top/processor/sha_core/n3636_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [1]),
	.I3(\top/processor/sha_core/w[57] [1]),
	.F(\top/processor/sha_core/n3637_170 )
);
defparam \top/processor/sha_core/n3637_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3496_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3868_131 ),
	.I3(\top/processor/sha_core/n3496_179 ),
	.F(\top/processor/sha_core/n3496_169 )
);
defparam \top/processor/sha_core/n3496_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3496_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [23]),
	.I2(\top/processor/sha_core/w[57] [23]),
	.F(\top/processor/sha_core/n3496_170 )
);
defparam \top/processor/sha_core/n3496_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [23]),
	.I2(\top/processor/sha_core/w[61] [23]),
	.F(\top/processor/sha_core/n3496_171 )
);
defparam \top/processor/sha_core/n3496_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3868_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3496_179 ),
	.I3(\top/processor/sha_core/n3496_170 ),
	.F(\top/processor/sha_core/n3868_130 )
);
defparam \top/processor/sha_core/n3868_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3868_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [23]),
	.I2(\top/processor/sha_core/w[63] [23]),
	.F(\top/processor/sha_core/n3868_131 )
);
defparam \top/processor/sha_core/n3868_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3638_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[59] [0]),
	.I3(\top/processor/sha_core/w[57] [0]),
	.F(\top/processor/sha_core/n3638_170 )
);
defparam \top/processor/sha_core/n3638_s149 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3497_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_117 ),
	.I3(\top/processor/sha_core/n3497_172 ),
	.F(\top/processor/sha_core/n3497_148 )
);
defparam \top/processor/sha_core/n3497_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [22]),
	.I2(\top/processor/sha_core/w[1] [22]),
	.F(\top/processor/sha_core/n3497_149 )
);
defparam \top/processor/sha_core/n3497_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [22]),
	.I2(\top/processor/sha_core/w[5] [22]),
	.F(\top/processor/sha_core/n3497_150 )
);
defparam \top/processor/sha_core/n3497_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_172 ),
	.I3(\top/processor/sha_core/n3497_149 ),
	.F(\top/processor/sha_core/n3869_116 )
);
defparam \top/processor/sha_core/n3869_s103 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3869_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [22]),
	.I2(\top/processor/sha_core/w[7] [22]),
	.F(\top/processor/sha_core/n3869_117 )
);
defparam \top/processor/sha_core/n3869_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [31]),
	.I3(\top/processor/sha_core/w[61] [31]),
	.F(\top/processor/sha_core/n3607_171 )
);
defparam \top/processor/sha_core/n3607_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [30]),
	.I3(\top/processor/sha_core/w[61] [30]),
	.F(\top/processor/sha_core/n3608_171 )
);
defparam \top/processor/sha_core/n3608_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [29]),
	.I3(\top/processor/sha_core/w[61] [29]),
	.F(\top/processor/sha_core/n3609_171 )
);
defparam \top/processor/sha_core/n3609_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [28]),
	.I3(\top/processor/sha_core/w[61] [28]),
	.F(\top/processor/sha_core/n3610_171 )
);
defparam \top/processor/sha_core/n3610_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [27]),
	.I3(\top/processor/sha_core/w[61] [27]),
	.F(\top/processor/sha_core/n3611_171 )
);
defparam \top/processor/sha_core/n3611_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [26]),
	.I3(\top/processor/sha_core/w[61] [26]),
	.F(\top/processor/sha_core/n3612_171 )
);
defparam \top/processor/sha_core/n3612_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [25]),
	.I3(\top/processor/sha_core/w[61] [25]),
	.F(\top/processor/sha_core/n3613_171 )
);
defparam \top/processor/sha_core/n3613_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3497_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_119 ),
	.I3(\top/processor/sha_core/n3497_173 ),
	.F(\top/processor/sha_core/n3497_151 )
);
defparam \top/processor/sha_core/n3497_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [22]),
	.I2(\top/processor/sha_core/w[9] [22]),
	.F(\top/processor/sha_core/n3497_152 )
);
defparam \top/processor/sha_core/n3497_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [22]),
	.I2(\top/processor/sha_core/w[13] [22]),
	.F(\top/processor/sha_core/n3497_153 )
);
defparam \top/processor/sha_core/n3497_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_173 ),
	.I3(\top/processor/sha_core/n3497_152 ),
	.F(\top/processor/sha_core/n3869_118 )
);
defparam \top/processor/sha_core/n3869_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [22]),
	.I2(\top/processor/sha_core/w[15] [22]),
	.F(\top/processor/sha_core/n3869_119 )
);
defparam \top/processor/sha_core/n3869_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3614_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [24]),
	.I3(\top/processor/sha_core/w[61] [24]),
	.F(\top/processor/sha_core/n3614_171 )
);
defparam \top/processor/sha_core/n3614_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [23]),
	.I3(\top/processor/sha_core/w[61] [23]),
	.F(\top/processor/sha_core/n3615_171 )
);
defparam \top/processor/sha_core/n3615_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [22]),
	.I3(\top/processor/sha_core/w[61] [22]),
	.F(\top/processor/sha_core/n3616_171 )
);
defparam \top/processor/sha_core/n3616_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [21]),
	.I3(\top/processor/sha_core/w[61] [21]),
	.F(\top/processor/sha_core/n3617_171 )
);
defparam \top/processor/sha_core/n3617_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [20]),
	.I3(\top/processor/sha_core/w[61] [20]),
	.F(\top/processor/sha_core/n3618_171 )
);
defparam \top/processor/sha_core/n3618_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [19]),
	.I3(\top/processor/sha_core/w[61] [19]),
	.F(\top/processor/sha_core/n3619_171 )
);
defparam \top/processor/sha_core/n3619_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [18]),
	.I3(\top/processor/sha_core/w[61] [18]),
	.F(\top/processor/sha_core/n3620_171 )
);
defparam \top/processor/sha_core/n3620_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [17]),
	.I3(\top/processor/sha_core/w[61] [17]),
	.F(\top/processor/sha_core/n3621_171 )
);
defparam \top/processor/sha_core/n3621_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [16]),
	.I3(\top/processor/sha_core/w[61] [16]),
	.F(\top/processor/sha_core/n3622_171 )
);
defparam \top/processor/sha_core/n3622_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [15]),
	.I3(\top/processor/sha_core/w[61] [15]),
	.F(\top/processor/sha_core/n3623_171 )
);
defparam \top/processor/sha_core/n3623_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [14]),
	.I3(\top/processor/sha_core/w[61] [14]),
	.F(\top/processor/sha_core/n3624_171 )
);
defparam \top/processor/sha_core/n3624_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [13]),
	.I3(\top/processor/sha_core/w[61] [13]),
	.F(\top/processor/sha_core/n3625_171 )
);
defparam \top/processor/sha_core/n3625_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [12]),
	.I3(\top/processor/sha_core/w[61] [12]),
	.F(\top/processor/sha_core/n3626_171 )
);
defparam \top/processor/sha_core/n3626_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [11]),
	.I3(\top/processor/sha_core/w[61] [11]),
	.F(\top/processor/sha_core/n3627_171 )
);
defparam \top/processor/sha_core/n3627_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [10]),
	.I3(\top/processor/sha_core/w[61] [10]),
	.F(\top/processor/sha_core/n3628_171 )
);
defparam \top/processor/sha_core/n3628_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [9]),
	.I3(\top/processor/sha_core/w[61] [9]),
	.F(\top/processor/sha_core/n3629_171 )
);
defparam \top/processor/sha_core/n3629_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [8]),
	.I3(\top/processor/sha_core/w[61] [8]),
	.F(\top/processor/sha_core/n3630_171 )
);
defparam \top/processor/sha_core/n3630_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [7]),
	.I3(\top/processor/sha_core/w[61] [7]),
	.F(\top/processor/sha_core/n3631_171 )
);
defparam \top/processor/sha_core/n3631_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [6]),
	.I3(\top/processor/sha_core/w[61] [6]),
	.F(\top/processor/sha_core/n3632_171 )
);
defparam \top/processor/sha_core/n3632_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [5]),
	.I3(\top/processor/sha_core/w[61] [5]),
	.F(\top/processor/sha_core/n3633_171 )
);
defparam \top/processor/sha_core/n3633_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3497_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_121 ),
	.I3(\top/processor/sha_core/n3497_174 ),
	.F(\top/processor/sha_core/n3497_154 )
);
defparam \top/processor/sha_core/n3497_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [22]),
	.I2(\top/processor/sha_core/w[17] [22]),
	.F(\top/processor/sha_core/n3497_155 )
);
defparam \top/processor/sha_core/n3497_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [22]),
	.I2(\top/processor/sha_core/w[21] [22]),
	.F(\top/processor/sha_core/n3497_156 )
);
defparam \top/processor/sha_core/n3497_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_174 ),
	.I3(\top/processor/sha_core/n3497_155 ),
	.F(\top/processor/sha_core/n3869_120 )
);
defparam \top/processor/sha_core/n3869_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [22]),
	.I2(\top/processor/sha_core/w[23] [22]),
	.F(\top/processor/sha_core/n3869_121 )
);
defparam \top/processor/sha_core/n3869_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3634_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [4]),
	.I3(\top/processor/sha_core/w[61] [4]),
	.F(\top/processor/sha_core/n3634_171 )
);
defparam \top/processor/sha_core/n3634_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [3]),
	.I3(\top/processor/sha_core/w[61] [3]),
	.F(\top/processor/sha_core/n3635_171 )
);
defparam \top/processor/sha_core/n3635_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [2]),
	.I3(\top/processor/sha_core/w[61] [2]),
	.F(\top/processor/sha_core/n3636_171 )
);
defparam \top/processor/sha_core/n3636_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [1]),
	.I3(\top/processor/sha_core/w[61] [1]),
	.F(\top/processor/sha_core/n3637_171 )
);
defparam \top/processor/sha_core/n3637_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s150  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[63] [0]),
	.I3(\top/processor/sha_core/w[61] [0]),
	.F(\top/processor/sha_core/n3638_171 )
);
defparam \top/processor/sha_core/n3638_s150 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3497_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_123 ),
	.I3(\top/processor/sha_core/n3497_175 ),
	.F(\top/processor/sha_core/n3497_157 )
);
defparam \top/processor/sha_core/n3497_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [22]),
	.I2(\top/processor/sha_core/w[25] [22]),
	.F(\top/processor/sha_core/n3497_158 )
);
defparam \top/processor/sha_core/n3497_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [22]),
	.I2(\top/processor/sha_core/w[29] [22]),
	.F(\top/processor/sha_core/n3497_159 )
);
defparam \top/processor/sha_core/n3497_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_175 ),
	.I3(\top/processor/sha_core/n3497_158 ),
	.F(\top/processor/sha_core/n3869_122 )
);
defparam \top/processor/sha_core/n3869_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [22]),
	.I2(\top/processor/sha_core/w[31] [22]),
	.F(\top/processor/sha_core/n3869_123 )
);
defparam \top/processor/sha_core/n3869_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3497_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_125 ),
	.I3(\top/processor/sha_core/n3497_176 ),
	.F(\top/processor/sha_core/n3497_160 )
);
defparam \top/processor/sha_core/n3497_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [22]),
	.I2(\top/processor/sha_core/w[33] [22]),
	.F(\top/processor/sha_core/n3497_161 )
);
defparam \top/processor/sha_core/n3497_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [22]),
	.I2(\top/processor/sha_core/w[37] [22]),
	.F(\top/processor/sha_core/n3497_162 )
);
defparam \top/processor/sha_core/n3497_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_176 ),
	.I3(\top/processor/sha_core/n3497_161 ),
	.F(\top/processor/sha_core/n3869_124 )
);
defparam \top/processor/sha_core/n3869_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [22]),
	.I2(\top/processor/sha_core/w[39] [22]),
	.F(\top/processor/sha_core/n3869_125 )
);
defparam \top/processor/sha_core/n3869_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3497_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_127 ),
	.I3(\top/processor/sha_core/n3497_177 ),
	.F(\top/processor/sha_core/n3497_163 )
);
defparam \top/processor/sha_core/n3497_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [22]),
	.I2(\top/processor/sha_core/w[41] [22]),
	.F(\top/processor/sha_core/n3497_164 )
);
defparam \top/processor/sha_core/n3497_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [22]),
	.I2(\top/processor/sha_core/w[45] [22]),
	.F(\top/processor/sha_core/n3497_165 )
);
defparam \top/processor/sha_core/n3497_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_177 ),
	.I3(\top/processor/sha_core/n3497_164 ),
	.F(\top/processor/sha_core/n3869_126 )
);
defparam \top/processor/sha_core/n3869_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [22]),
	.I2(\top/processor/sha_core/w[47] [22]),
	.F(\top/processor/sha_core/n3869_127 )
);
defparam \top/processor/sha_core/n3869_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3497_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_129 ),
	.I3(\top/processor/sha_core/n3497_178 ),
	.F(\top/processor/sha_core/n3497_166 )
);
defparam \top/processor/sha_core/n3497_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [22]),
	.I2(\top/processor/sha_core/w[49] [22]),
	.F(\top/processor/sha_core/n3497_167 )
);
defparam \top/processor/sha_core/n3497_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [22]),
	.I2(\top/processor/sha_core/w[53] [22]),
	.F(\top/processor/sha_core/n3497_168 )
);
defparam \top/processor/sha_core/n3497_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_178 ),
	.I3(\top/processor/sha_core/n3497_167 ),
	.F(\top/processor/sha_core/n3869_128 )
);
defparam \top/processor/sha_core/n3869_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [22]),
	.I2(\top/processor/sha_core/w[55] [22]),
	.F(\top/processor/sha_core/n3869_129 )
);
defparam \top/processor/sha_core/n3869_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3497_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3869_131 ),
	.I3(\top/processor/sha_core/n3497_179 ),
	.F(\top/processor/sha_core/n3497_169 )
);
defparam \top/processor/sha_core/n3497_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3497_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [22]),
	.I2(\top/processor/sha_core/w[57] [22]),
	.F(\top/processor/sha_core/n3497_170 )
);
defparam \top/processor/sha_core/n3497_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [22]),
	.I2(\top/processor/sha_core/w[61] [22]),
	.F(\top/processor/sha_core/n3497_171 )
);
defparam \top/processor/sha_core/n3497_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3869_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3497_179 ),
	.I3(\top/processor/sha_core/n3497_170 ),
	.F(\top/processor/sha_core/n3869_130 )
);
defparam \top/processor/sha_core/n3869_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3869_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [22]),
	.I2(\top/processor/sha_core/w[63] [22]),
	.F(\top/processor/sha_core/n3869_131 )
);
defparam \top/processor/sha_core/n3869_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_121 ),
	.I3(\top/processor/sha_core/n3488_174 ),
	.F(\top/processor/sha_core/n3488_154 )
);
defparam \top/processor/sha_core/n3488_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [31]),
	.I2(\top/processor/sha_core/w[57] [31]),
	.F(\top/processor/sha_core/n3488_155 )
);
defparam \top/processor/sha_core/n3488_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [31]),
	.I2(\top/processor/sha_core/w[61] [31]),
	.F(\top/processor/sha_core/n3488_156 )
);
defparam \top/processor/sha_core/n3488_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_174 ),
	.I3(\top/processor/sha_core/n3488_155 ),
	.F(\top/processor/sha_core/n3860_120 )
);
defparam \top/processor/sha_core/n3860_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [31]),
	.I2(\top/processor/sha_core/w[63] [31]),
	.F(\top/processor/sha_core/n3860_121 )
);
defparam \top/processor/sha_core/n3860_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_117 ),
	.I3(\top/processor/sha_core/n3498_172 ),
	.F(\top/processor/sha_core/n3498_148 )
);
defparam \top/processor/sha_core/n3498_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [21]),
	.I2(\top/processor/sha_core/w[1] [21]),
	.F(\top/processor/sha_core/n3498_149 )
);
defparam \top/processor/sha_core/n3498_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [21]),
	.I2(\top/processor/sha_core/w[5] [21]),
	.F(\top/processor/sha_core/n3498_150 )
);
defparam \top/processor/sha_core/n3498_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_172 ),
	.I3(\top/processor/sha_core/n3498_149 ),
	.F(\top/processor/sha_core/n3870_116 )
);
defparam \top/processor/sha_core/n3870_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [21]),
	.I2(\top/processor/sha_core/w[7] [21]),
	.F(\top/processor/sha_core/n3870_117 )
);
defparam \top/processor/sha_core/n3870_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_119 ),
	.I3(\top/processor/sha_core/n3498_173 ),
	.F(\top/processor/sha_core/n3498_151 )
);
defparam \top/processor/sha_core/n3498_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [21]),
	.I2(\top/processor/sha_core/w[9] [21]),
	.F(\top/processor/sha_core/n3498_152 )
);
defparam \top/processor/sha_core/n3498_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [21]),
	.I2(\top/processor/sha_core/w[13] [21]),
	.F(\top/processor/sha_core/n3498_153 )
);
defparam \top/processor/sha_core/n3498_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_173 ),
	.I3(\top/processor/sha_core/n3498_152 ),
	.F(\top/processor/sha_core/n3870_118 )
);
defparam \top/processor/sha_core/n3870_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [21]),
	.I2(\top/processor/sha_core/w[15] [21]),
	.F(\top/processor/sha_core/n3870_119 )
);
defparam \top/processor/sha_core/n3870_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_121 ),
	.I3(\top/processor/sha_core/n3498_174 ),
	.F(\top/processor/sha_core/n3498_154 )
);
defparam \top/processor/sha_core/n3498_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [21]),
	.I2(\top/processor/sha_core/w[17] [21]),
	.F(\top/processor/sha_core/n3498_155 )
);
defparam \top/processor/sha_core/n3498_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [21]),
	.I2(\top/processor/sha_core/w[21] [21]),
	.F(\top/processor/sha_core/n3498_156 )
);
defparam \top/processor/sha_core/n3498_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_174 ),
	.I3(\top/processor/sha_core/n3498_155 ),
	.F(\top/processor/sha_core/n3870_120 )
);
defparam \top/processor/sha_core/n3870_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [21]),
	.I2(\top/processor/sha_core/w[23] [21]),
	.F(\top/processor/sha_core/n3870_121 )
);
defparam \top/processor/sha_core/n3870_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_123 ),
	.I3(\top/processor/sha_core/n3498_175 ),
	.F(\top/processor/sha_core/n3498_157 )
);
defparam \top/processor/sha_core/n3498_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [21]),
	.I2(\top/processor/sha_core/w[25] [21]),
	.F(\top/processor/sha_core/n3498_158 )
);
defparam \top/processor/sha_core/n3498_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [21]),
	.I2(\top/processor/sha_core/w[29] [21]),
	.F(\top/processor/sha_core/n3498_159 )
);
defparam \top/processor/sha_core/n3498_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_175 ),
	.I3(\top/processor/sha_core/n3498_158 ),
	.F(\top/processor/sha_core/n3870_122 )
);
defparam \top/processor/sha_core/n3870_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [21]),
	.I2(\top/processor/sha_core/w[31] [21]),
	.F(\top/processor/sha_core/n3870_123 )
);
defparam \top/processor/sha_core/n3870_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_125 ),
	.I3(\top/processor/sha_core/n3498_176 ),
	.F(\top/processor/sha_core/n3498_160 )
);
defparam \top/processor/sha_core/n3498_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [21]),
	.I2(\top/processor/sha_core/w[33] [21]),
	.F(\top/processor/sha_core/n3498_161 )
);
defparam \top/processor/sha_core/n3498_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [21]),
	.I2(\top/processor/sha_core/w[37] [21]),
	.F(\top/processor/sha_core/n3498_162 )
);
defparam \top/processor/sha_core/n3498_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_176 ),
	.I3(\top/processor/sha_core/n3498_161 ),
	.F(\top/processor/sha_core/n3870_124 )
);
defparam \top/processor/sha_core/n3870_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [21]),
	.I2(\top/processor/sha_core/w[39] [21]),
	.F(\top/processor/sha_core/n3870_125 )
);
defparam \top/processor/sha_core/n3870_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_127 ),
	.I3(\top/processor/sha_core/n3498_177 ),
	.F(\top/processor/sha_core/n3498_163 )
);
defparam \top/processor/sha_core/n3498_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [21]),
	.I2(\top/processor/sha_core/w[41] [21]),
	.F(\top/processor/sha_core/n3498_164 )
);
defparam \top/processor/sha_core/n3498_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [21]),
	.I2(\top/processor/sha_core/w[45] [21]),
	.F(\top/processor/sha_core/n3498_165 )
);
defparam \top/processor/sha_core/n3498_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_177 ),
	.I3(\top/processor/sha_core/n3498_164 ),
	.F(\top/processor/sha_core/n3870_126 )
);
defparam \top/processor/sha_core/n3870_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [21]),
	.I2(\top/processor/sha_core/w[47] [21]),
	.F(\top/processor/sha_core/n3870_127 )
);
defparam \top/processor/sha_core/n3870_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_129 ),
	.I3(\top/processor/sha_core/n3498_178 ),
	.F(\top/processor/sha_core/n3498_166 )
);
defparam \top/processor/sha_core/n3498_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [21]),
	.I2(\top/processor/sha_core/w[49] [21]),
	.F(\top/processor/sha_core/n3498_167 )
);
defparam \top/processor/sha_core/n3498_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [21]),
	.I2(\top/processor/sha_core/w[53] [21]),
	.F(\top/processor/sha_core/n3498_168 )
);
defparam \top/processor/sha_core/n3498_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_178 ),
	.I3(\top/processor/sha_core/n3498_167 ),
	.F(\top/processor/sha_core/n3870_128 )
);
defparam \top/processor/sha_core/n3870_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [21]),
	.I2(\top/processor/sha_core/w[55] [21]),
	.F(\top/processor/sha_core/n3870_129 )
);
defparam \top/processor/sha_core/n3870_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3498_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3870_131 ),
	.I3(\top/processor/sha_core/n3498_179 ),
	.F(\top/processor/sha_core/n3498_169 )
);
defparam \top/processor/sha_core/n3498_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3498_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [21]),
	.I2(\top/processor/sha_core/w[57] [21]),
	.F(\top/processor/sha_core/n3498_170 )
);
defparam \top/processor/sha_core/n3498_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [21]),
	.I2(\top/processor/sha_core/w[61] [21]),
	.F(\top/processor/sha_core/n3498_171 )
);
defparam \top/processor/sha_core/n3498_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3870_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3498_179 ),
	.I3(\top/processor/sha_core/n3498_170 ),
	.F(\top/processor/sha_core/n3870_130 )
);
defparam \top/processor/sha_core/n3870_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3870_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [21]),
	.I2(\top/processor/sha_core/w[63] [21]),
	.F(\top/processor/sha_core/n3870_131 )
);
defparam \top/processor/sha_core/n3870_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_117 ),
	.I3(\top/processor/sha_core/n3499_172 ),
	.F(\top/processor/sha_core/n3499_148 )
);
defparam \top/processor/sha_core/n3499_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [20]),
	.I2(\top/processor/sha_core/w[1] [20]),
	.F(\top/processor/sha_core/n3499_149 )
);
defparam \top/processor/sha_core/n3499_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [20]),
	.I2(\top/processor/sha_core/w[5] [20]),
	.F(\top/processor/sha_core/n3499_150 )
);
defparam \top/processor/sha_core/n3499_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_172 ),
	.I3(\top/processor/sha_core/n3499_149 ),
	.F(\top/processor/sha_core/n3871_116 )
);
defparam \top/processor/sha_core/n3871_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [20]),
	.I2(\top/processor/sha_core/w[7] [20]),
	.F(\top/processor/sha_core/n3871_117 )
);
defparam \top/processor/sha_core/n3871_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_119 ),
	.I3(\top/processor/sha_core/n3499_173 ),
	.F(\top/processor/sha_core/n3499_151 )
);
defparam \top/processor/sha_core/n3499_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [20]),
	.I2(\top/processor/sha_core/w[9] [20]),
	.F(\top/processor/sha_core/n3499_152 )
);
defparam \top/processor/sha_core/n3499_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [20]),
	.I2(\top/processor/sha_core/w[13] [20]),
	.F(\top/processor/sha_core/n3499_153 )
);
defparam \top/processor/sha_core/n3499_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_173 ),
	.I3(\top/processor/sha_core/n3499_152 ),
	.F(\top/processor/sha_core/n3871_118 )
);
defparam \top/processor/sha_core/n3871_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [20]),
	.I2(\top/processor/sha_core/w[15] [20]),
	.F(\top/processor/sha_core/n3871_119 )
);
defparam \top/processor/sha_core/n3871_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_117 ),
	.I3(\top/processor/sha_core/n3489_172 ),
	.F(\top/processor/sha_core/n3489_148 )
);
defparam \top/processor/sha_core/n3489_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [30]),
	.I2(\top/processor/sha_core/w[1] [30]),
	.F(\top/processor/sha_core/n3489_149 )
);
defparam \top/processor/sha_core/n3489_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [30]),
	.I2(\top/processor/sha_core/w[5] [30]),
	.F(\top/processor/sha_core/n3489_150 )
);
defparam \top/processor/sha_core/n3489_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_172 ),
	.I3(\top/processor/sha_core/n3489_149 ),
	.F(\top/processor/sha_core/n3861_116 )
);
defparam \top/processor/sha_core/n3861_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [30]),
	.I2(\top/processor/sha_core/w[7] [30]),
	.F(\top/processor/sha_core/n3861_117 )
);
defparam \top/processor/sha_core/n3861_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_121 ),
	.I3(\top/processor/sha_core/n3499_174 ),
	.F(\top/processor/sha_core/n3499_154 )
);
defparam \top/processor/sha_core/n3499_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [20]),
	.I2(\top/processor/sha_core/w[17] [20]),
	.F(\top/processor/sha_core/n3499_155 )
);
defparam \top/processor/sha_core/n3499_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [20]),
	.I2(\top/processor/sha_core/w[21] [20]),
	.F(\top/processor/sha_core/n3499_156 )
);
defparam \top/processor/sha_core/n3499_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_174 ),
	.I3(\top/processor/sha_core/n3499_155 ),
	.F(\top/processor/sha_core/n3871_120 )
);
defparam \top/processor/sha_core/n3871_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [20]),
	.I2(\top/processor/sha_core/w[23] [20]),
	.F(\top/processor/sha_core/n3871_121 )
);
defparam \top/processor/sha_core/n3871_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_123 ),
	.I3(\top/processor/sha_core/n3499_175 ),
	.F(\top/processor/sha_core/n3499_157 )
);
defparam \top/processor/sha_core/n3499_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [20]),
	.I2(\top/processor/sha_core/w[25] [20]),
	.F(\top/processor/sha_core/n3499_158 )
);
defparam \top/processor/sha_core/n3499_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [20]),
	.I2(\top/processor/sha_core/w[29] [20]),
	.F(\top/processor/sha_core/n3499_159 )
);
defparam \top/processor/sha_core/n3499_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_175 ),
	.I3(\top/processor/sha_core/n3499_158 ),
	.F(\top/processor/sha_core/n3871_122 )
);
defparam \top/processor/sha_core/n3871_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [20]),
	.I2(\top/processor/sha_core/w[31] [20]),
	.F(\top/processor/sha_core/n3871_123 )
);
defparam \top/processor/sha_core/n3871_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_125 ),
	.I3(\top/processor/sha_core/n3499_176 ),
	.F(\top/processor/sha_core/n3499_160 )
);
defparam \top/processor/sha_core/n3499_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [20]),
	.I2(\top/processor/sha_core/w[33] [20]),
	.F(\top/processor/sha_core/n3499_161 )
);
defparam \top/processor/sha_core/n3499_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [20]),
	.I2(\top/processor/sha_core/w[37] [20]),
	.F(\top/processor/sha_core/n3499_162 )
);
defparam \top/processor/sha_core/n3499_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_176 ),
	.I3(\top/processor/sha_core/n3499_161 ),
	.F(\top/processor/sha_core/n3871_124 )
);
defparam \top/processor/sha_core/n3871_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [20]),
	.I2(\top/processor/sha_core/w[39] [20]),
	.F(\top/processor/sha_core/n3871_125 )
);
defparam \top/processor/sha_core/n3871_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_127 ),
	.I3(\top/processor/sha_core/n3499_177 ),
	.F(\top/processor/sha_core/n3499_163 )
);
defparam \top/processor/sha_core/n3499_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [20]),
	.I2(\top/processor/sha_core/w[41] [20]),
	.F(\top/processor/sha_core/n3499_164 )
);
defparam \top/processor/sha_core/n3499_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [20]),
	.I2(\top/processor/sha_core/w[45] [20]),
	.F(\top/processor/sha_core/n3499_165 )
);
defparam \top/processor/sha_core/n3499_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_177 ),
	.I3(\top/processor/sha_core/n3499_164 ),
	.F(\top/processor/sha_core/n3871_126 )
);
defparam \top/processor/sha_core/n3871_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [20]),
	.I2(\top/processor/sha_core/w[47] [20]),
	.F(\top/processor/sha_core/n3871_127 )
);
defparam \top/processor/sha_core/n3871_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_129 ),
	.I3(\top/processor/sha_core/n3499_178 ),
	.F(\top/processor/sha_core/n3499_166 )
);
defparam \top/processor/sha_core/n3499_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [20]),
	.I2(\top/processor/sha_core/w[49] [20]),
	.F(\top/processor/sha_core/n3499_167 )
);
defparam \top/processor/sha_core/n3499_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [20]),
	.I2(\top/processor/sha_core/w[53] [20]),
	.F(\top/processor/sha_core/n3499_168 )
);
defparam \top/processor/sha_core/n3499_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_178 ),
	.I3(\top/processor/sha_core/n3499_167 ),
	.F(\top/processor/sha_core/n3871_128 )
);
defparam \top/processor/sha_core/n3871_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [20]),
	.I2(\top/processor/sha_core/w[55] [20]),
	.F(\top/processor/sha_core/n3871_129 )
);
defparam \top/processor/sha_core/n3871_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3499_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3871_131 ),
	.I3(\top/processor/sha_core/n3499_179 ),
	.F(\top/processor/sha_core/n3499_169 )
);
defparam \top/processor/sha_core/n3499_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3499_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [20]),
	.I2(\top/processor/sha_core/w[57] [20]),
	.F(\top/processor/sha_core/n3499_170 )
);
defparam \top/processor/sha_core/n3499_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [20]),
	.I2(\top/processor/sha_core/w[61] [20]),
	.F(\top/processor/sha_core/n3499_171 )
);
defparam \top/processor/sha_core/n3499_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3871_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3499_179 ),
	.I3(\top/processor/sha_core/n3499_170 ),
	.F(\top/processor/sha_core/n3871_130 )
);
defparam \top/processor/sha_core/n3871_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3871_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [20]),
	.I2(\top/processor/sha_core/w[63] [20]),
	.F(\top/processor/sha_core/n3871_131 )
);
defparam \top/processor/sha_core/n3871_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_117 ),
	.I3(\top/processor/sha_core/n3500_172 ),
	.F(\top/processor/sha_core/n3500_148 )
);
defparam \top/processor/sha_core/n3500_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [19]),
	.I2(\top/processor/sha_core/w[1] [19]),
	.F(\top/processor/sha_core/n3500_149 )
);
defparam \top/processor/sha_core/n3500_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [19]),
	.I2(\top/processor/sha_core/w[5] [19]),
	.F(\top/processor/sha_core/n3500_150 )
);
defparam \top/processor/sha_core/n3500_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_172 ),
	.I3(\top/processor/sha_core/n3500_149 ),
	.F(\top/processor/sha_core/n3872_116 )
);
defparam \top/processor/sha_core/n3872_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [19]),
	.I2(\top/processor/sha_core/w[7] [19]),
	.F(\top/processor/sha_core/n3872_117 )
);
defparam \top/processor/sha_core/n3872_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_119 ),
	.I3(\top/processor/sha_core/n3500_173 ),
	.F(\top/processor/sha_core/n3500_151 )
);
defparam \top/processor/sha_core/n3500_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [19]),
	.I2(\top/processor/sha_core/w[9] [19]),
	.F(\top/processor/sha_core/n3500_152 )
);
defparam \top/processor/sha_core/n3500_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [19]),
	.I2(\top/processor/sha_core/w[13] [19]),
	.F(\top/processor/sha_core/n3500_153 )
);
defparam \top/processor/sha_core/n3500_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_173 ),
	.I3(\top/processor/sha_core/n3500_152 ),
	.F(\top/processor/sha_core/n3872_118 )
);
defparam \top/processor/sha_core/n3872_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [19]),
	.I2(\top/processor/sha_core/w[15] [19]),
	.F(\top/processor/sha_core/n3872_119 )
);
defparam \top/processor/sha_core/n3872_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_121 ),
	.I3(\top/processor/sha_core/n3500_174 ),
	.F(\top/processor/sha_core/n3500_154 )
);
defparam \top/processor/sha_core/n3500_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [19]),
	.I2(\top/processor/sha_core/w[17] [19]),
	.F(\top/processor/sha_core/n3500_155 )
);
defparam \top/processor/sha_core/n3500_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [19]),
	.I2(\top/processor/sha_core/w[21] [19]),
	.F(\top/processor/sha_core/n3500_156 )
);
defparam \top/processor/sha_core/n3500_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_174 ),
	.I3(\top/processor/sha_core/n3500_155 ),
	.F(\top/processor/sha_core/n3872_120 )
);
defparam \top/processor/sha_core/n3872_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [19]),
	.I2(\top/processor/sha_core/w[23] [19]),
	.F(\top/processor/sha_core/n3872_121 )
);
defparam \top/processor/sha_core/n3872_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_123 ),
	.I3(\top/processor/sha_core/n3500_175 ),
	.F(\top/processor/sha_core/n3500_157 )
);
defparam \top/processor/sha_core/n3500_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [19]),
	.I2(\top/processor/sha_core/w[25] [19]),
	.F(\top/processor/sha_core/n3500_158 )
);
defparam \top/processor/sha_core/n3500_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [19]),
	.I2(\top/processor/sha_core/w[29] [19]),
	.F(\top/processor/sha_core/n3500_159 )
);
defparam \top/processor/sha_core/n3500_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_175 ),
	.I3(\top/processor/sha_core/n3500_158 ),
	.F(\top/processor/sha_core/n3872_122 )
);
defparam \top/processor/sha_core/n3872_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [19]),
	.I2(\top/processor/sha_core/w[31] [19]),
	.F(\top/processor/sha_core/n3872_123 )
);
defparam \top/processor/sha_core/n3872_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_119 ),
	.I3(\top/processor/sha_core/n3489_173 ),
	.F(\top/processor/sha_core/n3489_151 )
);
defparam \top/processor/sha_core/n3489_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [30]),
	.I2(\top/processor/sha_core/w[9] [30]),
	.F(\top/processor/sha_core/n3489_152 )
);
defparam \top/processor/sha_core/n3489_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [30]),
	.I2(\top/processor/sha_core/w[13] [30]),
	.F(\top/processor/sha_core/n3489_153 )
);
defparam \top/processor/sha_core/n3489_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_173 ),
	.I3(\top/processor/sha_core/n3489_152 ),
	.F(\top/processor/sha_core/n3861_118 )
);
defparam \top/processor/sha_core/n3861_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [30]),
	.I2(\top/processor/sha_core/w[15] [30]),
	.F(\top/processor/sha_core/n3861_119 )
);
defparam \top/processor/sha_core/n3861_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_123 ),
	.I3(\top/processor/sha_core/n3488_175 ),
	.F(\top/processor/sha_core/n3488_157 )
);
defparam \top/processor/sha_core/n3488_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [31]),
	.I2(\top/processor/sha_core/w[1] [31]),
	.F(\top/processor/sha_core/n3488_158 )
);
defparam \top/processor/sha_core/n3488_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [31]),
	.I2(\top/processor/sha_core/w[5] [31]),
	.F(\top/processor/sha_core/n3488_159 )
);
defparam \top/processor/sha_core/n3488_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_175 ),
	.I3(\top/processor/sha_core/n3488_158 ),
	.F(\top/processor/sha_core/n3860_122 )
);
defparam \top/processor/sha_core/n3860_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [31]),
	.I2(\top/processor/sha_core/w[7] [31]),
	.F(\top/processor/sha_core/n3860_123 )
);
defparam \top/processor/sha_core/n3860_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_125 ),
	.I3(\top/processor/sha_core/n3500_176 ),
	.F(\top/processor/sha_core/n3500_160 )
);
defparam \top/processor/sha_core/n3500_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [19]),
	.I2(\top/processor/sha_core/w[33] [19]),
	.F(\top/processor/sha_core/n3500_161 )
);
defparam \top/processor/sha_core/n3500_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [19]),
	.I2(\top/processor/sha_core/w[37] [19]),
	.F(\top/processor/sha_core/n3500_162 )
);
defparam \top/processor/sha_core/n3500_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_176 ),
	.I3(\top/processor/sha_core/n3500_161 ),
	.F(\top/processor/sha_core/n3872_124 )
);
defparam \top/processor/sha_core/n3872_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [19]),
	.I2(\top/processor/sha_core/w[39] [19]),
	.F(\top/processor/sha_core/n3872_125 )
);
defparam \top/processor/sha_core/n3872_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_127 ),
	.I3(\top/processor/sha_core/n3500_177 ),
	.F(\top/processor/sha_core/n3500_163 )
);
defparam \top/processor/sha_core/n3500_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [19]),
	.I2(\top/processor/sha_core/w[41] [19]),
	.F(\top/processor/sha_core/n3500_164 )
);
defparam \top/processor/sha_core/n3500_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [19]),
	.I2(\top/processor/sha_core/w[45] [19]),
	.F(\top/processor/sha_core/n3500_165 )
);
defparam \top/processor/sha_core/n3500_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_177 ),
	.I3(\top/processor/sha_core/n3500_164 ),
	.F(\top/processor/sha_core/n3872_126 )
);
defparam \top/processor/sha_core/n3872_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [19]),
	.I2(\top/processor/sha_core/w[47] [19]),
	.F(\top/processor/sha_core/n3872_127 )
);
defparam \top/processor/sha_core/n3872_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_129 ),
	.I3(\top/processor/sha_core/n3500_178 ),
	.F(\top/processor/sha_core/n3500_166 )
);
defparam \top/processor/sha_core/n3500_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [19]),
	.I2(\top/processor/sha_core/w[49] [19]),
	.F(\top/processor/sha_core/n3500_167 )
);
defparam \top/processor/sha_core/n3500_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [19]),
	.I2(\top/processor/sha_core/w[53] [19]),
	.F(\top/processor/sha_core/n3500_168 )
);
defparam \top/processor/sha_core/n3500_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_178 ),
	.I3(\top/processor/sha_core/n3500_167 ),
	.F(\top/processor/sha_core/n3872_128 )
);
defparam \top/processor/sha_core/n3872_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [19]),
	.I2(\top/processor/sha_core/w[55] [19]),
	.F(\top/processor/sha_core/n3872_129 )
);
defparam \top/processor/sha_core/n3872_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3500_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3872_131 ),
	.I3(\top/processor/sha_core/n3500_179 ),
	.F(\top/processor/sha_core/n3500_169 )
);
defparam \top/processor/sha_core/n3500_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3500_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [19]),
	.I2(\top/processor/sha_core/w[57] [19]),
	.F(\top/processor/sha_core/n3500_170 )
);
defparam \top/processor/sha_core/n3500_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [19]),
	.I2(\top/processor/sha_core/w[61] [19]),
	.F(\top/processor/sha_core/n3500_171 )
);
defparam \top/processor/sha_core/n3500_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3872_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3500_179 ),
	.I3(\top/processor/sha_core/n3500_170 ),
	.F(\top/processor/sha_core/n3872_130 )
);
defparam \top/processor/sha_core/n3872_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3872_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [19]),
	.I2(\top/processor/sha_core/w[63] [19]),
	.F(\top/processor/sha_core/n3872_131 )
);
defparam \top/processor/sha_core/n3872_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_117 ),
	.I3(\top/processor/sha_core/n3501_172 ),
	.F(\top/processor/sha_core/n3501_148 )
);
defparam \top/processor/sha_core/n3501_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [18]),
	.I2(\top/processor/sha_core/w[1] [18]),
	.F(\top/processor/sha_core/n3501_149 )
);
defparam \top/processor/sha_core/n3501_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [18]),
	.I2(\top/processor/sha_core/w[5] [18]),
	.F(\top/processor/sha_core/n3501_150 )
);
defparam \top/processor/sha_core/n3501_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_172 ),
	.I3(\top/processor/sha_core/n3501_149 ),
	.F(\top/processor/sha_core/n3873_116 )
);
defparam \top/processor/sha_core/n3873_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [18]),
	.I2(\top/processor/sha_core/w[7] [18]),
	.F(\top/processor/sha_core/n3873_117 )
);
defparam \top/processor/sha_core/n3873_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_119 ),
	.I3(\top/processor/sha_core/n3501_173 ),
	.F(\top/processor/sha_core/n3501_151 )
);
defparam \top/processor/sha_core/n3501_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [18]),
	.I2(\top/processor/sha_core/w[9] [18]),
	.F(\top/processor/sha_core/n3501_152 )
);
defparam \top/processor/sha_core/n3501_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [18]),
	.I2(\top/processor/sha_core/w[13] [18]),
	.F(\top/processor/sha_core/n3501_153 )
);
defparam \top/processor/sha_core/n3501_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_173 ),
	.I3(\top/processor/sha_core/n3501_152 ),
	.F(\top/processor/sha_core/n3873_118 )
);
defparam \top/processor/sha_core/n3873_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [18]),
	.I2(\top/processor/sha_core/w[15] [18]),
	.F(\top/processor/sha_core/n3873_119 )
);
defparam \top/processor/sha_core/n3873_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_121 ),
	.I3(\top/processor/sha_core/n3501_174 ),
	.F(\top/processor/sha_core/n3501_154 )
);
defparam \top/processor/sha_core/n3501_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [18]),
	.I2(\top/processor/sha_core/w[17] [18]),
	.F(\top/processor/sha_core/n3501_155 )
);
defparam \top/processor/sha_core/n3501_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [18]),
	.I2(\top/processor/sha_core/w[21] [18]),
	.F(\top/processor/sha_core/n3501_156 )
);
defparam \top/processor/sha_core/n3501_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_174 ),
	.I3(\top/processor/sha_core/n3501_155 ),
	.F(\top/processor/sha_core/n3873_120 )
);
defparam \top/processor/sha_core/n3873_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [18]),
	.I2(\top/processor/sha_core/w[23] [18]),
	.F(\top/processor/sha_core/n3873_121 )
);
defparam \top/processor/sha_core/n3873_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_123 ),
	.I3(\top/processor/sha_core/n3501_175 ),
	.F(\top/processor/sha_core/n3501_157 )
);
defparam \top/processor/sha_core/n3501_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [18]),
	.I2(\top/processor/sha_core/w[25] [18]),
	.F(\top/processor/sha_core/n3501_158 )
);
defparam \top/processor/sha_core/n3501_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [18]),
	.I2(\top/processor/sha_core/w[29] [18]),
	.F(\top/processor/sha_core/n3501_159 )
);
defparam \top/processor/sha_core/n3501_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_175 ),
	.I3(\top/processor/sha_core/n3501_158 ),
	.F(\top/processor/sha_core/n3873_122 )
);
defparam \top/processor/sha_core/n3873_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [18]),
	.I2(\top/processor/sha_core/w[31] [18]),
	.F(\top/processor/sha_core/n3873_123 )
);
defparam \top/processor/sha_core/n3873_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_125 ),
	.I3(\top/processor/sha_core/n3501_176 ),
	.F(\top/processor/sha_core/n3501_160 )
);
defparam \top/processor/sha_core/n3501_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [18]),
	.I2(\top/processor/sha_core/w[33] [18]),
	.F(\top/processor/sha_core/n3501_161 )
);
defparam \top/processor/sha_core/n3501_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [18]),
	.I2(\top/processor/sha_core/w[37] [18]),
	.F(\top/processor/sha_core/n3501_162 )
);
defparam \top/processor/sha_core/n3501_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_176 ),
	.I3(\top/processor/sha_core/n3501_161 ),
	.F(\top/processor/sha_core/n3873_124 )
);
defparam \top/processor/sha_core/n3873_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [18]),
	.I2(\top/processor/sha_core/w[39] [18]),
	.F(\top/processor/sha_core/n3873_125 )
);
defparam \top/processor/sha_core/n3873_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_127 ),
	.I3(\top/processor/sha_core/n3501_177 ),
	.F(\top/processor/sha_core/n3501_163 )
);
defparam \top/processor/sha_core/n3501_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [18]),
	.I2(\top/processor/sha_core/w[41] [18]),
	.F(\top/processor/sha_core/n3501_164 )
);
defparam \top/processor/sha_core/n3501_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [18]),
	.I2(\top/processor/sha_core/w[45] [18]),
	.F(\top/processor/sha_core/n3501_165 )
);
defparam \top/processor/sha_core/n3501_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_177 ),
	.I3(\top/processor/sha_core/n3501_164 ),
	.F(\top/processor/sha_core/n3873_126 )
);
defparam \top/processor/sha_core/n3873_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [18]),
	.I2(\top/processor/sha_core/w[47] [18]),
	.F(\top/processor/sha_core/n3873_127 )
);
defparam \top/processor/sha_core/n3873_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_121 ),
	.I3(\top/processor/sha_core/n3489_174 ),
	.F(\top/processor/sha_core/n3489_154 )
);
defparam \top/processor/sha_core/n3489_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [30]),
	.I2(\top/processor/sha_core/w[17] [30]),
	.F(\top/processor/sha_core/n3489_155 )
);
defparam \top/processor/sha_core/n3489_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [30]),
	.I2(\top/processor/sha_core/w[21] [30]),
	.F(\top/processor/sha_core/n3489_156 )
);
defparam \top/processor/sha_core/n3489_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_174 ),
	.I3(\top/processor/sha_core/n3489_155 ),
	.F(\top/processor/sha_core/n3861_120 )
);
defparam \top/processor/sha_core/n3861_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [30]),
	.I2(\top/processor/sha_core/w[23] [30]),
	.F(\top/processor/sha_core/n3861_121 )
);
defparam \top/processor/sha_core/n3861_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_129 ),
	.I3(\top/processor/sha_core/n3501_178 ),
	.F(\top/processor/sha_core/n3501_166 )
);
defparam \top/processor/sha_core/n3501_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [18]),
	.I2(\top/processor/sha_core/w[49] [18]),
	.F(\top/processor/sha_core/n3501_167 )
);
defparam \top/processor/sha_core/n3501_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [18]),
	.I2(\top/processor/sha_core/w[53] [18]),
	.F(\top/processor/sha_core/n3501_168 )
);
defparam \top/processor/sha_core/n3501_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_178 ),
	.I3(\top/processor/sha_core/n3501_167 ),
	.F(\top/processor/sha_core/n3873_128 )
);
defparam \top/processor/sha_core/n3873_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [18]),
	.I2(\top/processor/sha_core/w[55] [18]),
	.F(\top/processor/sha_core/n3873_129 )
);
defparam \top/processor/sha_core/n3873_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3501_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3873_131 ),
	.I3(\top/processor/sha_core/n3501_179 ),
	.F(\top/processor/sha_core/n3501_169 )
);
defparam \top/processor/sha_core/n3501_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3501_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [18]),
	.I2(\top/processor/sha_core/w[57] [18]),
	.F(\top/processor/sha_core/n3501_170 )
);
defparam \top/processor/sha_core/n3501_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [18]),
	.I2(\top/processor/sha_core/w[61] [18]),
	.F(\top/processor/sha_core/n3501_171 )
);
defparam \top/processor/sha_core/n3501_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3873_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3501_179 ),
	.I3(\top/processor/sha_core/n3501_170 ),
	.F(\top/processor/sha_core/n3873_130 )
);
defparam \top/processor/sha_core/n3873_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3873_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [18]),
	.I2(\top/processor/sha_core/w[63] [18]),
	.F(\top/processor/sha_core/n3873_131 )
);
defparam \top/processor/sha_core/n3873_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_117 ),
	.I3(\top/processor/sha_core/n3502_172 ),
	.F(\top/processor/sha_core/n3502_148 )
);
defparam \top/processor/sha_core/n3502_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [17]),
	.I2(\top/processor/sha_core/w[1] [17]),
	.F(\top/processor/sha_core/n3502_149 )
);
defparam \top/processor/sha_core/n3502_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [17]),
	.I2(\top/processor/sha_core/w[5] [17]),
	.F(\top/processor/sha_core/n3502_150 )
);
defparam \top/processor/sha_core/n3502_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_172 ),
	.I3(\top/processor/sha_core/n3502_149 ),
	.F(\top/processor/sha_core/n3874_116 )
);
defparam \top/processor/sha_core/n3874_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [17]),
	.I2(\top/processor/sha_core/w[7] [17]),
	.F(\top/processor/sha_core/n3874_117 )
);
defparam \top/processor/sha_core/n3874_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_119 ),
	.I3(\top/processor/sha_core/n3502_173 ),
	.F(\top/processor/sha_core/n3502_151 )
);
defparam \top/processor/sha_core/n3502_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [17]),
	.I2(\top/processor/sha_core/w[9] [17]),
	.F(\top/processor/sha_core/n3502_152 )
);
defparam \top/processor/sha_core/n3502_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [17]),
	.I2(\top/processor/sha_core/w[13] [17]),
	.F(\top/processor/sha_core/n3502_153 )
);
defparam \top/processor/sha_core/n3502_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_173 ),
	.I3(\top/processor/sha_core/n3502_152 ),
	.F(\top/processor/sha_core/n3874_118 )
);
defparam \top/processor/sha_core/n3874_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [17]),
	.I2(\top/processor/sha_core/w[15] [17]),
	.F(\top/processor/sha_core/n3874_119 )
);
defparam \top/processor/sha_core/n3874_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_121 ),
	.I3(\top/processor/sha_core/n3502_174 ),
	.F(\top/processor/sha_core/n3502_154 )
);
defparam \top/processor/sha_core/n3502_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [17]),
	.I2(\top/processor/sha_core/w[17] [17]),
	.F(\top/processor/sha_core/n3502_155 )
);
defparam \top/processor/sha_core/n3502_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [17]),
	.I2(\top/processor/sha_core/w[21] [17]),
	.F(\top/processor/sha_core/n3502_156 )
);
defparam \top/processor/sha_core/n3502_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_174 ),
	.I3(\top/processor/sha_core/n3502_155 ),
	.F(\top/processor/sha_core/n3874_120 )
);
defparam \top/processor/sha_core/n3874_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [17]),
	.I2(\top/processor/sha_core/w[23] [17]),
	.F(\top/processor/sha_core/n3874_121 )
);
defparam \top/processor/sha_core/n3874_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_123 ),
	.I3(\top/processor/sha_core/n3502_175 ),
	.F(\top/processor/sha_core/n3502_157 )
);
defparam \top/processor/sha_core/n3502_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [17]),
	.I2(\top/processor/sha_core/w[25] [17]),
	.F(\top/processor/sha_core/n3502_158 )
);
defparam \top/processor/sha_core/n3502_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [17]),
	.I2(\top/processor/sha_core/w[29] [17]),
	.F(\top/processor/sha_core/n3502_159 )
);
defparam \top/processor/sha_core/n3502_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_175 ),
	.I3(\top/processor/sha_core/n3502_158 ),
	.F(\top/processor/sha_core/n3874_122 )
);
defparam \top/processor/sha_core/n3874_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [17]),
	.I2(\top/processor/sha_core/w[31] [17]),
	.F(\top/processor/sha_core/n3874_123 )
);
defparam \top/processor/sha_core/n3874_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_125 ),
	.I3(\top/processor/sha_core/n3502_176 ),
	.F(\top/processor/sha_core/n3502_160 )
);
defparam \top/processor/sha_core/n3502_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [17]),
	.I2(\top/processor/sha_core/w[33] [17]),
	.F(\top/processor/sha_core/n3502_161 )
);
defparam \top/processor/sha_core/n3502_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [17]),
	.I2(\top/processor/sha_core/w[37] [17]),
	.F(\top/processor/sha_core/n3502_162 )
);
defparam \top/processor/sha_core/n3502_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_176 ),
	.I3(\top/processor/sha_core/n3502_161 ),
	.F(\top/processor/sha_core/n3874_124 )
);
defparam \top/processor/sha_core/n3874_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [17]),
	.I2(\top/processor/sha_core/w[39] [17]),
	.F(\top/processor/sha_core/n3874_125 )
);
defparam \top/processor/sha_core/n3874_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_127 ),
	.I3(\top/processor/sha_core/n3502_177 ),
	.F(\top/processor/sha_core/n3502_163 )
);
defparam \top/processor/sha_core/n3502_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [17]),
	.I2(\top/processor/sha_core/w[41] [17]),
	.F(\top/processor/sha_core/n3502_164 )
);
defparam \top/processor/sha_core/n3502_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [17]),
	.I2(\top/processor/sha_core/w[45] [17]),
	.F(\top/processor/sha_core/n3502_165 )
);
defparam \top/processor/sha_core/n3502_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_177 ),
	.I3(\top/processor/sha_core/n3502_164 ),
	.F(\top/processor/sha_core/n3874_126 )
);
defparam \top/processor/sha_core/n3874_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [17]),
	.I2(\top/processor/sha_core/w[47] [17]),
	.F(\top/processor/sha_core/n3874_127 )
);
defparam \top/processor/sha_core/n3874_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_129 ),
	.I3(\top/processor/sha_core/n3502_178 ),
	.F(\top/processor/sha_core/n3502_166 )
);
defparam \top/processor/sha_core/n3502_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [17]),
	.I2(\top/processor/sha_core/w[49] [17]),
	.F(\top/processor/sha_core/n3502_167 )
);
defparam \top/processor/sha_core/n3502_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [17]),
	.I2(\top/processor/sha_core/w[53] [17]),
	.F(\top/processor/sha_core/n3502_168 )
);
defparam \top/processor/sha_core/n3502_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_178 ),
	.I3(\top/processor/sha_core/n3502_167 ),
	.F(\top/processor/sha_core/n3874_128 )
);
defparam \top/processor/sha_core/n3874_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [17]),
	.I2(\top/processor/sha_core/w[55] [17]),
	.F(\top/processor/sha_core/n3874_129 )
);
defparam \top/processor/sha_core/n3874_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3502_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3874_131 ),
	.I3(\top/processor/sha_core/n3502_179 ),
	.F(\top/processor/sha_core/n3502_169 )
);
defparam \top/processor/sha_core/n3502_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3502_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [17]),
	.I2(\top/processor/sha_core/w[57] [17]),
	.F(\top/processor/sha_core/n3502_170 )
);
defparam \top/processor/sha_core/n3502_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [17]),
	.I2(\top/processor/sha_core/w[61] [17]),
	.F(\top/processor/sha_core/n3502_171 )
);
defparam \top/processor/sha_core/n3502_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3874_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3502_179 ),
	.I3(\top/processor/sha_core/n3502_170 ),
	.F(\top/processor/sha_core/n3874_130 )
);
defparam \top/processor/sha_core/n3874_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3874_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [17]),
	.I2(\top/processor/sha_core/w[63] [17]),
	.F(\top/processor/sha_core/n3874_131 )
);
defparam \top/processor/sha_core/n3874_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_123 ),
	.I3(\top/processor/sha_core/n3489_175 ),
	.F(\top/processor/sha_core/n3489_157 )
);
defparam \top/processor/sha_core/n3489_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [30]),
	.I2(\top/processor/sha_core/w[25] [30]),
	.F(\top/processor/sha_core/n3489_158 )
);
defparam \top/processor/sha_core/n3489_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [30]),
	.I2(\top/processor/sha_core/w[29] [30]),
	.F(\top/processor/sha_core/n3489_159 )
);
defparam \top/processor/sha_core/n3489_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_175 ),
	.I3(\top/processor/sha_core/n3489_158 ),
	.F(\top/processor/sha_core/n3861_122 )
);
defparam \top/processor/sha_core/n3861_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [30]),
	.I2(\top/processor/sha_core/w[31] [30]),
	.F(\top/processor/sha_core/n3861_123 )
);
defparam \top/processor/sha_core/n3861_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_117 ),
	.I3(\top/processor/sha_core/n3503_172 ),
	.F(\top/processor/sha_core/n3503_148 )
);
defparam \top/processor/sha_core/n3503_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [16]),
	.I2(\top/processor/sha_core/w[1] [16]),
	.F(\top/processor/sha_core/n3503_149 )
);
defparam \top/processor/sha_core/n3503_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [16]),
	.I2(\top/processor/sha_core/w[5] [16]),
	.F(\top/processor/sha_core/n3503_150 )
);
defparam \top/processor/sha_core/n3503_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_172 ),
	.I3(\top/processor/sha_core/n3503_149 ),
	.F(\top/processor/sha_core/n3875_116 )
);
defparam \top/processor/sha_core/n3875_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [16]),
	.I2(\top/processor/sha_core/w[7] [16]),
	.F(\top/processor/sha_core/n3875_117 )
);
defparam \top/processor/sha_core/n3875_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_119 ),
	.I3(\top/processor/sha_core/n3503_173 ),
	.F(\top/processor/sha_core/n3503_151 )
);
defparam \top/processor/sha_core/n3503_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [16]),
	.I2(\top/processor/sha_core/w[9] [16]),
	.F(\top/processor/sha_core/n3503_152 )
);
defparam \top/processor/sha_core/n3503_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [16]),
	.I2(\top/processor/sha_core/w[13] [16]),
	.F(\top/processor/sha_core/n3503_153 )
);
defparam \top/processor/sha_core/n3503_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_173 ),
	.I3(\top/processor/sha_core/n3503_152 ),
	.F(\top/processor/sha_core/n3875_118 )
);
defparam \top/processor/sha_core/n3875_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [16]),
	.I2(\top/processor/sha_core/w[15] [16]),
	.F(\top/processor/sha_core/n3875_119 )
);
defparam \top/processor/sha_core/n3875_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_121 ),
	.I3(\top/processor/sha_core/n3503_174 ),
	.F(\top/processor/sha_core/n3503_154 )
);
defparam \top/processor/sha_core/n3503_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [16]),
	.I2(\top/processor/sha_core/w[17] [16]),
	.F(\top/processor/sha_core/n3503_155 )
);
defparam \top/processor/sha_core/n3503_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [16]),
	.I2(\top/processor/sha_core/w[21] [16]),
	.F(\top/processor/sha_core/n3503_156 )
);
defparam \top/processor/sha_core/n3503_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_174 ),
	.I3(\top/processor/sha_core/n3503_155 ),
	.F(\top/processor/sha_core/n3875_120 )
);
defparam \top/processor/sha_core/n3875_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [16]),
	.I2(\top/processor/sha_core/w[23] [16]),
	.F(\top/processor/sha_core/n3875_121 )
);
defparam \top/processor/sha_core/n3875_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_123 ),
	.I3(\top/processor/sha_core/n3503_175 ),
	.F(\top/processor/sha_core/n3503_157 )
);
defparam \top/processor/sha_core/n3503_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [16]),
	.I2(\top/processor/sha_core/w[25] [16]),
	.F(\top/processor/sha_core/n3503_158 )
);
defparam \top/processor/sha_core/n3503_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [16]),
	.I2(\top/processor/sha_core/w[29] [16]),
	.F(\top/processor/sha_core/n3503_159 )
);
defparam \top/processor/sha_core/n3503_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_175 ),
	.I3(\top/processor/sha_core/n3503_158 ),
	.F(\top/processor/sha_core/n3875_122 )
);
defparam \top/processor/sha_core/n3875_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [16]),
	.I2(\top/processor/sha_core/w[31] [16]),
	.F(\top/processor/sha_core/n3875_123 )
);
defparam \top/processor/sha_core/n3875_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_125 ),
	.I3(\top/processor/sha_core/n3503_176 ),
	.F(\top/processor/sha_core/n3503_160 )
);
defparam \top/processor/sha_core/n3503_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [16]),
	.I2(\top/processor/sha_core/w[33] [16]),
	.F(\top/processor/sha_core/n3503_161 )
);
defparam \top/processor/sha_core/n3503_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [16]),
	.I2(\top/processor/sha_core/w[37] [16]),
	.F(\top/processor/sha_core/n3503_162 )
);
defparam \top/processor/sha_core/n3503_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_176 ),
	.I3(\top/processor/sha_core/n3503_161 ),
	.F(\top/processor/sha_core/n3875_124 )
);
defparam \top/processor/sha_core/n3875_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [16]),
	.I2(\top/processor/sha_core/w[39] [16]),
	.F(\top/processor/sha_core/n3875_125 )
);
defparam \top/processor/sha_core/n3875_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_127 ),
	.I3(\top/processor/sha_core/n3503_177 ),
	.F(\top/processor/sha_core/n3503_163 )
);
defparam \top/processor/sha_core/n3503_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [16]),
	.I2(\top/processor/sha_core/w[41] [16]),
	.F(\top/processor/sha_core/n3503_164 )
);
defparam \top/processor/sha_core/n3503_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [16]),
	.I2(\top/processor/sha_core/w[45] [16]),
	.F(\top/processor/sha_core/n3503_165 )
);
defparam \top/processor/sha_core/n3503_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_177 ),
	.I3(\top/processor/sha_core/n3503_164 ),
	.F(\top/processor/sha_core/n3875_126 )
);
defparam \top/processor/sha_core/n3875_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [16]),
	.I2(\top/processor/sha_core/w[47] [16]),
	.F(\top/processor/sha_core/n3875_127 )
);
defparam \top/processor/sha_core/n3875_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_129 ),
	.I3(\top/processor/sha_core/n3503_178 ),
	.F(\top/processor/sha_core/n3503_166 )
);
defparam \top/processor/sha_core/n3503_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [16]),
	.I2(\top/processor/sha_core/w[49] [16]),
	.F(\top/processor/sha_core/n3503_167 )
);
defparam \top/processor/sha_core/n3503_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [16]),
	.I2(\top/processor/sha_core/w[53] [16]),
	.F(\top/processor/sha_core/n3503_168 )
);
defparam \top/processor/sha_core/n3503_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_178 ),
	.I3(\top/processor/sha_core/n3503_167 ),
	.F(\top/processor/sha_core/n3875_128 )
);
defparam \top/processor/sha_core/n3875_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [16]),
	.I2(\top/processor/sha_core/w[55] [16]),
	.F(\top/processor/sha_core/n3875_129 )
);
defparam \top/processor/sha_core/n3875_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3503_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3875_131 ),
	.I3(\top/processor/sha_core/n3503_179 ),
	.F(\top/processor/sha_core/n3503_169 )
);
defparam \top/processor/sha_core/n3503_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3503_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [16]),
	.I2(\top/processor/sha_core/w[57] [16]),
	.F(\top/processor/sha_core/n3503_170 )
);
defparam \top/processor/sha_core/n3503_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [16]),
	.I2(\top/processor/sha_core/w[61] [16]),
	.F(\top/processor/sha_core/n3503_171 )
);
defparam \top/processor/sha_core/n3503_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3875_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3503_179 ),
	.I3(\top/processor/sha_core/n3503_170 ),
	.F(\top/processor/sha_core/n3875_130 )
);
defparam \top/processor/sha_core/n3875_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3875_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [16]),
	.I2(\top/processor/sha_core/w[63] [16]),
	.F(\top/processor/sha_core/n3875_131 )
);
defparam \top/processor/sha_core/n3875_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_117 ),
	.I3(\top/processor/sha_core/n3504_172 ),
	.F(\top/processor/sha_core/n3504_148 )
);
defparam \top/processor/sha_core/n3504_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [15]),
	.I2(\top/processor/sha_core/w[1] [15]),
	.F(\top/processor/sha_core/n3504_149 )
);
defparam \top/processor/sha_core/n3504_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [15]),
	.I2(\top/processor/sha_core/w[5] [15]),
	.F(\top/processor/sha_core/n3504_150 )
);
defparam \top/processor/sha_core/n3504_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_172 ),
	.I3(\top/processor/sha_core/n3504_149 ),
	.F(\top/processor/sha_core/n3876_116 )
);
defparam \top/processor/sha_core/n3876_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [15]),
	.I2(\top/processor/sha_core/w[7] [15]),
	.F(\top/processor/sha_core/n3876_117 )
);
defparam \top/processor/sha_core/n3876_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_119 ),
	.I3(\top/processor/sha_core/n3504_173 ),
	.F(\top/processor/sha_core/n3504_151 )
);
defparam \top/processor/sha_core/n3504_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [15]),
	.I2(\top/processor/sha_core/w[9] [15]),
	.F(\top/processor/sha_core/n3504_152 )
);
defparam \top/processor/sha_core/n3504_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [15]),
	.I2(\top/processor/sha_core/w[13] [15]),
	.F(\top/processor/sha_core/n3504_153 )
);
defparam \top/processor/sha_core/n3504_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_173 ),
	.I3(\top/processor/sha_core/n3504_152 ),
	.F(\top/processor/sha_core/n3876_118 )
);
defparam \top/processor/sha_core/n3876_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [15]),
	.I2(\top/processor/sha_core/w[15] [15]),
	.F(\top/processor/sha_core/n3876_119 )
);
defparam \top/processor/sha_core/n3876_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_125 ),
	.I3(\top/processor/sha_core/n3489_176 ),
	.F(\top/processor/sha_core/n3489_160 )
);
defparam \top/processor/sha_core/n3489_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [30]),
	.I2(\top/processor/sha_core/w[33] [30]),
	.F(\top/processor/sha_core/n3489_161 )
);
defparam \top/processor/sha_core/n3489_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [30]),
	.I2(\top/processor/sha_core/w[37] [30]),
	.F(\top/processor/sha_core/n3489_162 )
);
defparam \top/processor/sha_core/n3489_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_176 ),
	.I3(\top/processor/sha_core/n3489_161 ),
	.F(\top/processor/sha_core/n3861_124 )
);
defparam \top/processor/sha_core/n3861_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [30]),
	.I2(\top/processor/sha_core/w[39] [30]),
	.F(\top/processor/sha_core/n3861_125 )
);
defparam \top/processor/sha_core/n3861_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_121 ),
	.I3(\top/processor/sha_core/n3504_174 ),
	.F(\top/processor/sha_core/n3504_154 )
);
defparam \top/processor/sha_core/n3504_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [15]),
	.I2(\top/processor/sha_core/w[17] [15]),
	.F(\top/processor/sha_core/n3504_155 )
);
defparam \top/processor/sha_core/n3504_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [15]),
	.I2(\top/processor/sha_core/w[21] [15]),
	.F(\top/processor/sha_core/n3504_156 )
);
defparam \top/processor/sha_core/n3504_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_174 ),
	.I3(\top/processor/sha_core/n3504_155 ),
	.F(\top/processor/sha_core/n3876_120 )
);
defparam \top/processor/sha_core/n3876_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [15]),
	.I2(\top/processor/sha_core/w[23] [15]),
	.F(\top/processor/sha_core/n3876_121 )
);
defparam \top/processor/sha_core/n3876_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_123 ),
	.I3(\top/processor/sha_core/n3504_175 ),
	.F(\top/processor/sha_core/n3504_157 )
);
defparam \top/processor/sha_core/n3504_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [15]),
	.I2(\top/processor/sha_core/w[25] [15]),
	.F(\top/processor/sha_core/n3504_158 )
);
defparam \top/processor/sha_core/n3504_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [15]),
	.I2(\top/processor/sha_core/w[29] [15]),
	.F(\top/processor/sha_core/n3504_159 )
);
defparam \top/processor/sha_core/n3504_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_175 ),
	.I3(\top/processor/sha_core/n3504_158 ),
	.F(\top/processor/sha_core/n3876_122 )
);
defparam \top/processor/sha_core/n3876_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [15]),
	.I2(\top/processor/sha_core/w[31] [15]),
	.F(\top/processor/sha_core/n3876_123 )
);
defparam \top/processor/sha_core/n3876_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_125 ),
	.I3(\top/processor/sha_core/n3504_176 ),
	.F(\top/processor/sha_core/n3504_160 )
);
defparam \top/processor/sha_core/n3504_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [15]),
	.I2(\top/processor/sha_core/w[33] [15]),
	.F(\top/processor/sha_core/n3504_161 )
);
defparam \top/processor/sha_core/n3504_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [15]),
	.I2(\top/processor/sha_core/w[37] [15]),
	.F(\top/processor/sha_core/n3504_162 )
);
defparam \top/processor/sha_core/n3504_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_176 ),
	.I3(\top/processor/sha_core/n3504_161 ),
	.F(\top/processor/sha_core/n3876_124 )
);
defparam \top/processor/sha_core/n3876_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [15]),
	.I2(\top/processor/sha_core/w[39] [15]),
	.F(\top/processor/sha_core/n3876_125 )
);
defparam \top/processor/sha_core/n3876_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_127 ),
	.I3(\top/processor/sha_core/n3504_177 ),
	.F(\top/processor/sha_core/n3504_163 )
);
defparam \top/processor/sha_core/n3504_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [15]),
	.I2(\top/processor/sha_core/w[41] [15]),
	.F(\top/processor/sha_core/n3504_164 )
);
defparam \top/processor/sha_core/n3504_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [15]),
	.I2(\top/processor/sha_core/w[45] [15]),
	.F(\top/processor/sha_core/n3504_165 )
);
defparam \top/processor/sha_core/n3504_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_177 ),
	.I3(\top/processor/sha_core/n3504_164 ),
	.F(\top/processor/sha_core/n3876_126 )
);
defparam \top/processor/sha_core/n3876_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [15]),
	.I2(\top/processor/sha_core/w[47] [15]),
	.F(\top/processor/sha_core/n3876_127 )
);
defparam \top/processor/sha_core/n3876_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_129 ),
	.I3(\top/processor/sha_core/n3504_178 ),
	.F(\top/processor/sha_core/n3504_166 )
);
defparam \top/processor/sha_core/n3504_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [15]),
	.I2(\top/processor/sha_core/w[49] [15]),
	.F(\top/processor/sha_core/n3504_167 )
);
defparam \top/processor/sha_core/n3504_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [15]),
	.I2(\top/processor/sha_core/w[53] [15]),
	.F(\top/processor/sha_core/n3504_168 )
);
defparam \top/processor/sha_core/n3504_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_178 ),
	.I3(\top/processor/sha_core/n3504_167 ),
	.F(\top/processor/sha_core/n3876_128 )
);
defparam \top/processor/sha_core/n3876_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [15]),
	.I2(\top/processor/sha_core/w[55] [15]),
	.F(\top/processor/sha_core/n3876_129 )
);
defparam \top/processor/sha_core/n3876_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3504_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3876_131 ),
	.I3(\top/processor/sha_core/n3504_179 ),
	.F(\top/processor/sha_core/n3504_169 )
);
defparam \top/processor/sha_core/n3504_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3504_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [15]),
	.I2(\top/processor/sha_core/w[57] [15]),
	.F(\top/processor/sha_core/n3504_170 )
);
defparam \top/processor/sha_core/n3504_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [15]),
	.I2(\top/processor/sha_core/w[61] [15]),
	.F(\top/processor/sha_core/n3504_171 )
);
defparam \top/processor/sha_core/n3504_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3876_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3504_179 ),
	.I3(\top/processor/sha_core/n3504_170 ),
	.F(\top/processor/sha_core/n3876_130 )
);
defparam \top/processor/sha_core/n3876_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3876_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [15]),
	.I2(\top/processor/sha_core/w[63] [15]),
	.F(\top/processor/sha_core/n3876_131 )
);
defparam \top/processor/sha_core/n3876_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_117 ),
	.I3(\top/processor/sha_core/n3505_172 ),
	.F(\top/processor/sha_core/n3505_148 )
);
defparam \top/processor/sha_core/n3505_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [14]),
	.I2(\top/processor/sha_core/w[1] [14]),
	.F(\top/processor/sha_core/n3505_149 )
);
defparam \top/processor/sha_core/n3505_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [14]),
	.I2(\top/processor/sha_core/w[5] [14]),
	.F(\top/processor/sha_core/n3505_150 )
);
defparam \top/processor/sha_core/n3505_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_172 ),
	.I3(\top/processor/sha_core/n3505_149 ),
	.F(\top/processor/sha_core/n3877_116 )
);
defparam \top/processor/sha_core/n3877_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [14]),
	.I2(\top/processor/sha_core/w[7] [14]),
	.F(\top/processor/sha_core/n3877_117 )
);
defparam \top/processor/sha_core/n3877_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_119 ),
	.I3(\top/processor/sha_core/n3505_173 ),
	.F(\top/processor/sha_core/n3505_151 )
);
defparam \top/processor/sha_core/n3505_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [14]),
	.I2(\top/processor/sha_core/w[9] [14]),
	.F(\top/processor/sha_core/n3505_152 )
);
defparam \top/processor/sha_core/n3505_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [14]),
	.I2(\top/processor/sha_core/w[13] [14]),
	.F(\top/processor/sha_core/n3505_153 )
);
defparam \top/processor/sha_core/n3505_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_173 ),
	.I3(\top/processor/sha_core/n3505_152 ),
	.F(\top/processor/sha_core/n3877_118 )
);
defparam \top/processor/sha_core/n3877_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [14]),
	.I2(\top/processor/sha_core/w[15] [14]),
	.F(\top/processor/sha_core/n3877_119 )
);
defparam \top/processor/sha_core/n3877_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_121 ),
	.I3(\top/processor/sha_core/n3505_174 ),
	.F(\top/processor/sha_core/n3505_154 )
);
defparam \top/processor/sha_core/n3505_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [14]),
	.I2(\top/processor/sha_core/w[17] [14]),
	.F(\top/processor/sha_core/n3505_155 )
);
defparam \top/processor/sha_core/n3505_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [14]),
	.I2(\top/processor/sha_core/w[21] [14]),
	.F(\top/processor/sha_core/n3505_156 )
);
defparam \top/processor/sha_core/n3505_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_174 ),
	.I3(\top/processor/sha_core/n3505_155 ),
	.F(\top/processor/sha_core/n3877_120 )
);
defparam \top/processor/sha_core/n3877_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [14]),
	.I2(\top/processor/sha_core/w[23] [14]),
	.F(\top/processor/sha_core/n3877_121 )
);
defparam \top/processor/sha_core/n3877_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_123 ),
	.I3(\top/processor/sha_core/n3505_175 ),
	.F(\top/processor/sha_core/n3505_157 )
);
defparam \top/processor/sha_core/n3505_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [14]),
	.I2(\top/processor/sha_core/w[25] [14]),
	.F(\top/processor/sha_core/n3505_158 )
);
defparam \top/processor/sha_core/n3505_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [14]),
	.I2(\top/processor/sha_core/w[29] [14]),
	.F(\top/processor/sha_core/n3505_159 )
);
defparam \top/processor/sha_core/n3505_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_175 ),
	.I3(\top/processor/sha_core/n3505_158 ),
	.F(\top/processor/sha_core/n3877_122 )
);
defparam \top/processor/sha_core/n3877_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [14]),
	.I2(\top/processor/sha_core/w[31] [14]),
	.F(\top/processor/sha_core/n3877_123 )
);
defparam \top/processor/sha_core/n3877_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_127 ),
	.I3(\top/processor/sha_core/n3489_177 ),
	.F(\top/processor/sha_core/n3489_163 )
);
defparam \top/processor/sha_core/n3489_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [30]),
	.I2(\top/processor/sha_core/w[41] [30]),
	.F(\top/processor/sha_core/n3489_164 )
);
defparam \top/processor/sha_core/n3489_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [30]),
	.I2(\top/processor/sha_core/w[45] [30]),
	.F(\top/processor/sha_core/n3489_165 )
);
defparam \top/processor/sha_core/n3489_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_177 ),
	.I3(\top/processor/sha_core/n3489_164 ),
	.F(\top/processor/sha_core/n3861_126 )
);
defparam \top/processor/sha_core/n3861_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [30]),
	.I2(\top/processor/sha_core/w[47] [30]),
	.F(\top/processor/sha_core/n3861_127 )
);
defparam \top/processor/sha_core/n3861_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_125 ),
	.I3(\top/processor/sha_core/n3505_176 ),
	.F(\top/processor/sha_core/n3505_160 )
);
defparam \top/processor/sha_core/n3505_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [14]),
	.I2(\top/processor/sha_core/w[33] [14]),
	.F(\top/processor/sha_core/n3505_161 )
);
defparam \top/processor/sha_core/n3505_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [14]),
	.I2(\top/processor/sha_core/w[37] [14]),
	.F(\top/processor/sha_core/n3505_162 )
);
defparam \top/processor/sha_core/n3505_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_176 ),
	.I3(\top/processor/sha_core/n3505_161 ),
	.F(\top/processor/sha_core/n3877_124 )
);
defparam \top/processor/sha_core/n3877_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [14]),
	.I2(\top/processor/sha_core/w[39] [14]),
	.F(\top/processor/sha_core/n3877_125 )
);
defparam \top/processor/sha_core/n3877_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_127 ),
	.I3(\top/processor/sha_core/n3505_177 ),
	.F(\top/processor/sha_core/n3505_163 )
);
defparam \top/processor/sha_core/n3505_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [14]),
	.I2(\top/processor/sha_core/w[41] [14]),
	.F(\top/processor/sha_core/n3505_164 )
);
defparam \top/processor/sha_core/n3505_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [14]),
	.I2(\top/processor/sha_core/w[45] [14]),
	.F(\top/processor/sha_core/n3505_165 )
);
defparam \top/processor/sha_core/n3505_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_177 ),
	.I3(\top/processor/sha_core/n3505_164 ),
	.F(\top/processor/sha_core/n3877_126 )
);
defparam \top/processor/sha_core/n3877_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [14]),
	.I2(\top/processor/sha_core/w[47] [14]),
	.F(\top/processor/sha_core/n3877_127 )
);
defparam \top/processor/sha_core/n3877_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_129 ),
	.I3(\top/processor/sha_core/n3505_178 ),
	.F(\top/processor/sha_core/n3505_166 )
);
defparam \top/processor/sha_core/n3505_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [14]),
	.I2(\top/processor/sha_core/w[49] [14]),
	.F(\top/processor/sha_core/n3505_167 )
);
defparam \top/processor/sha_core/n3505_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [14]),
	.I2(\top/processor/sha_core/w[53] [14]),
	.F(\top/processor/sha_core/n3505_168 )
);
defparam \top/processor/sha_core/n3505_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_178 ),
	.I3(\top/processor/sha_core/n3505_167 ),
	.F(\top/processor/sha_core/n3877_128 )
);
defparam \top/processor/sha_core/n3877_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [14]),
	.I2(\top/processor/sha_core/w[55] [14]),
	.F(\top/processor/sha_core/n3877_129 )
);
defparam \top/processor/sha_core/n3877_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3505_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3877_131 ),
	.I3(\top/processor/sha_core/n3505_179 ),
	.F(\top/processor/sha_core/n3505_169 )
);
defparam \top/processor/sha_core/n3505_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3505_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [14]),
	.I2(\top/processor/sha_core/w[57] [14]),
	.F(\top/processor/sha_core/n3505_170 )
);
defparam \top/processor/sha_core/n3505_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [14]),
	.I2(\top/processor/sha_core/w[61] [14]),
	.F(\top/processor/sha_core/n3505_171 )
);
defparam \top/processor/sha_core/n3505_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3877_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3505_179 ),
	.I3(\top/processor/sha_core/n3505_170 ),
	.F(\top/processor/sha_core/n3877_130 )
);
defparam \top/processor/sha_core/n3877_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3877_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [14]),
	.I2(\top/processor/sha_core/w[63] [14]),
	.F(\top/processor/sha_core/n3877_131 )
);
defparam \top/processor/sha_core/n3877_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_117 ),
	.I3(\top/processor/sha_core/n3506_172 ),
	.F(\top/processor/sha_core/n3506_148 )
);
defparam \top/processor/sha_core/n3506_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [13]),
	.I2(\top/processor/sha_core/w[1] [13]),
	.F(\top/processor/sha_core/n3506_149 )
);
defparam \top/processor/sha_core/n3506_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [13]),
	.I2(\top/processor/sha_core/w[5] [13]),
	.F(\top/processor/sha_core/n3506_150 )
);
defparam \top/processor/sha_core/n3506_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_172 ),
	.I3(\top/processor/sha_core/n3506_149 ),
	.F(\top/processor/sha_core/n3878_116 )
);
defparam \top/processor/sha_core/n3878_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [13]),
	.I2(\top/processor/sha_core/w[7] [13]),
	.F(\top/processor/sha_core/n3878_117 )
);
defparam \top/processor/sha_core/n3878_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_119 ),
	.I3(\top/processor/sha_core/n3506_173 ),
	.F(\top/processor/sha_core/n3506_151 )
);
defparam \top/processor/sha_core/n3506_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [13]),
	.I2(\top/processor/sha_core/w[9] [13]),
	.F(\top/processor/sha_core/n3506_152 )
);
defparam \top/processor/sha_core/n3506_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [13]),
	.I2(\top/processor/sha_core/w[13] [13]),
	.F(\top/processor/sha_core/n3506_153 )
);
defparam \top/processor/sha_core/n3506_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_173 ),
	.I3(\top/processor/sha_core/n3506_152 ),
	.F(\top/processor/sha_core/n3878_118 )
);
defparam \top/processor/sha_core/n3878_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [13]),
	.I2(\top/processor/sha_core/w[15] [13]),
	.F(\top/processor/sha_core/n3878_119 )
);
defparam \top/processor/sha_core/n3878_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_121 ),
	.I3(\top/processor/sha_core/n3506_174 ),
	.F(\top/processor/sha_core/n3506_154 )
);
defparam \top/processor/sha_core/n3506_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [13]),
	.I2(\top/processor/sha_core/w[17] [13]),
	.F(\top/processor/sha_core/n3506_155 )
);
defparam \top/processor/sha_core/n3506_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [13]),
	.I2(\top/processor/sha_core/w[21] [13]),
	.F(\top/processor/sha_core/n3506_156 )
);
defparam \top/processor/sha_core/n3506_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_174 ),
	.I3(\top/processor/sha_core/n3506_155 ),
	.F(\top/processor/sha_core/n3878_120 )
);
defparam \top/processor/sha_core/n3878_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [13]),
	.I2(\top/processor/sha_core/w[23] [13]),
	.F(\top/processor/sha_core/n3878_121 )
);
defparam \top/processor/sha_core/n3878_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_123 ),
	.I3(\top/processor/sha_core/n3506_175 ),
	.F(\top/processor/sha_core/n3506_157 )
);
defparam \top/processor/sha_core/n3506_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [13]),
	.I2(\top/processor/sha_core/w[25] [13]),
	.F(\top/processor/sha_core/n3506_158 )
);
defparam \top/processor/sha_core/n3506_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [13]),
	.I2(\top/processor/sha_core/w[29] [13]),
	.F(\top/processor/sha_core/n3506_159 )
);
defparam \top/processor/sha_core/n3506_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_175 ),
	.I3(\top/processor/sha_core/n3506_158 ),
	.F(\top/processor/sha_core/n3878_122 )
);
defparam \top/processor/sha_core/n3878_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [13]),
	.I2(\top/processor/sha_core/w[31] [13]),
	.F(\top/processor/sha_core/n3878_123 )
);
defparam \top/processor/sha_core/n3878_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_125 ),
	.I3(\top/processor/sha_core/n3506_176 ),
	.F(\top/processor/sha_core/n3506_160 )
);
defparam \top/processor/sha_core/n3506_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [13]),
	.I2(\top/processor/sha_core/w[33] [13]),
	.F(\top/processor/sha_core/n3506_161 )
);
defparam \top/processor/sha_core/n3506_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [13]),
	.I2(\top/processor/sha_core/w[37] [13]),
	.F(\top/processor/sha_core/n3506_162 )
);
defparam \top/processor/sha_core/n3506_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_176 ),
	.I3(\top/processor/sha_core/n3506_161 ),
	.F(\top/processor/sha_core/n3878_124 )
);
defparam \top/processor/sha_core/n3878_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [13]),
	.I2(\top/processor/sha_core/w[39] [13]),
	.F(\top/processor/sha_core/n3878_125 )
);
defparam \top/processor/sha_core/n3878_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_127 ),
	.I3(\top/processor/sha_core/n3506_177 ),
	.F(\top/processor/sha_core/n3506_163 )
);
defparam \top/processor/sha_core/n3506_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [13]),
	.I2(\top/processor/sha_core/w[41] [13]),
	.F(\top/processor/sha_core/n3506_164 )
);
defparam \top/processor/sha_core/n3506_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [13]),
	.I2(\top/processor/sha_core/w[45] [13]),
	.F(\top/processor/sha_core/n3506_165 )
);
defparam \top/processor/sha_core/n3506_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_177 ),
	.I3(\top/processor/sha_core/n3506_164 ),
	.F(\top/processor/sha_core/n3878_126 )
);
defparam \top/processor/sha_core/n3878_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [13]),
	.I2(\top/processor/sha_core/w[47] [13]),
	.F(\top/processor/sha_core/n3878_127 )
);
defparam \top/processor/sha_core/n3878_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_129 ),
	.I3(\top/processor/sha_core/n3489_178 ),
	.F(\top/processor/sha_core/n3489_166 )
);
defparam \top/processor/sha_core/n3489_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [30]),
	.I2(\top/processor/sha_core/w[49] [30]),
	.F(\top/processor/sha_core/n3489_167 )
);
defparam \top/processor/sha_core/n3489_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [30]),
	.I2(\top/processor/sha_core/w[53] [30]),
	.F(\top/processor/sha_core/n3489_168 )
);
defparam \top/processor/sha_core/n3489_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_178 ),
	.I3(\top/processor/sha_core/n3489_167 ),
	.F(\top/processor/sha_core/n3861_128 )
);
defparam \top/processor/sha_core/n3861_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [30]),
	.I2(\top/processor/sha_core/w[55] [30]),
	.F(\top/processor/sha_core/n3861_129 )
);
defparam \top/processor/sha_core/n3861_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_129 ),
	.I3(\top/processor/sha_core/n3506_178 ),
	.F(\top/processor/sha_core/n3506_166 )
);
defparam \top/processor/sha_core/n3506_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [13]),
	.I2(\top/processor/sha_core/w[49] [13]),
	.F(\top/processor/sha_core/n3506_167 )
);
defparam \top/processor/sha_core/n3506_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [13]),
	.I2(\top/processor/sha_core/w[53] [13]),
	.F(\top/processor/sha_core/n3506_168 )
);
defparam \top/processor/sha_core/n3506_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_178 ),
	.I3(\top/processor/sha_core/n3506_167 ),
	.F(\top/processor/sha_core/n3878_128 )
);
defparam \top/processor/sha_core/n3878_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [13]),
	.I2(\top/processor/sha_core/w[55] [13]),
	.F(\top/processor/sha_core/n3878_129 )
);
defparam \top/processor/sha_core/n3878_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3506_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3878_131 ),
	.I3(\top/processor/sha_core/n3506_179 ),
	.F(\top/processor/sha_core/n3506_169 )
);
defparam \top/processor/sha_core/n3506_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3506_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [13]),
	.I2(\top/processor/sha_core/w[57] [13]),
	.F(\top/processor/sha_core/n3506_170 )
);
defparam \top/processor/sha_core/n3506_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [13]),
	.I2(\top/processor/sha_core/w[61] [13]),
	.F(\top/processor/sha_core/n3506_171 )
);
defparam \top/processor/sha_core/n3506_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3878_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3506_179 ),
	.I3(\top/processor/sha_core/n3506_170 ),
	.F(\top/processor/sha_core/n3878_130 )
);
defparam \top/processor/sha_core/n3878_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3878_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [13]),
	.I2(\top/processor/sha_core/w[63] [13]),
	.F(\top/processor/sha_core/n3878_131 )
);
defparam \top/processor/sha_core/n3878_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_117 ),
	.I3(\top/processor/sha_core/n3507_172 ),
	.F(\top/processor/sha_core/n3507_148 )
);
defparam \top/processor/sha_core/n3507_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [12]),
	.I2(\top/processor/sha_core/w[1] [12]),
	.F(\top/processor/sha_core/n3507_149 )
);
defparam \top/processor/sha_core/n3507_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [12]),
	.I2(\top/processor/sha_core/w[5] [12]),
	.F(\top/processor/sha_core/n3507_150 )
);
defparam \top/processor/sha_core/n3507_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_172 ),
	.I3(\top/processor/sha_core/n3507_149 ),
	.F(\top/processor/sha_core/n3879_116 )
);
defparam \top/processor/sha_core/n3879_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [12]),
	.I2(\top/processor/sha_core/w[7] [12]),
	.F(\top/processor/sha_core/n3879_117 )
);
defparam \top/processor/sha_core/n3879_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_119 ),
	.I3(\top/processor/sha_core/n3507_173 ),
	.F(\top/processor/sha_core/n3507_151 )
);
defparam \top/processor/sha_core/n3507_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [12]),
	.I2(\top/processor/sha_core/w[9] [12]),
	.F(\top/processor/sha_core/n3507_152 )
);
defparam \top/processor/sha_core/n3507_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [12]),
	.I2(\top/processor/sha_core/w[13] [12]),
	.F(\top/processor/sha_core/n3507_153 )
);
defparam \top/processor/sha_core/n3507_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_173 ),
	.I3(\top/processor/sha_core/n3507_152 ),
	.F(\top/processor/sha_core/n3879_118 )
);
defparam \top/processor/sha_core/n3879_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [12]),
	.I2(\top/processor/sha_core/w[15] [12]),
	.F(\top/processor/sha_core/n3879_119 )
);
defparam \top/processor/sha_core/n3879_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_121 ),
	.I3(\top/processor/sha_core/n3507_174 ),
	.F(\top/processor/sha_core/n3507_154 )
);
defparam \top/processor/sha_core/n3507_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [12]),
	.I2(\top/processor/sha_core/w[17] [12]),
	.F(\top/processor/sha_core/n3507_155 )
);
defparam \top/processor/sha_core/n3507_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [12]),
	.I2(\top/processor/sha_core/w[21] [12]),
	.F(\top/processor/sha_core/n3507_156 )
);
defparam \top/processor/sha_core/n3507_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_174 ),
	.I3(\top/processor/sha_core/n3507_155 ),
	.F(\top/processor/sha_core/n3879_120 )
);
defparam \top/processor/sha_core/n3879_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [12]),
	.I2(\top/processor/sha_core/w[23] [12]),
	.F(\top/processor/sha_core/n3879_121 )
);
defparam \top/processor/sha_core/n3879_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_123 ),
	.I3(\top/processor/sha_core/n3507_175 ),
	.F(\top/processor/sha_core/n3507_157 )
);
defparam \top/processor/sha_core/n3507_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [12]),
	.I2(\top/processor/sha_core/w[25] [12]),
	.F(\top/processor/sha_core/n3507_158 )
);
defparam \top/processor/sha_core/n3507_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [12]),
	.I2(\top/processor/sha_core/w[29] [12]),
	.F(\top/processor/sha_core/n3507_159 )
);
defparam \top/processor/sha_core/n3507_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_175 ),
	.I3(\top/processor/sha_core/n3507_158 ),
	.F(\top/processor/sha_core/n3879_122 )
);
defparam \top/processor/sha_core/n3879_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [12]),
	.I2(\top/processor/sha_core/w[31] [12]),
	.F(\top/processor/sha_core/n3879_123 )
);
defparam \top/processor/sha_core/n3879_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_125 ),
	.I3(\top/processor/sha_core/n3507_176 ),
	.F(\top/processor/sha_core/n3507_160 )
);
defparam \top/processor/sha_core/n3507_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [12]),
	.I2(\top/processor/sha_core/w[33] [12]),
	.F(\top/processor/sha_core/n3507_161 )
);
defparam \top/processor/sha_core/n3507_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [12]),
	.I2(\top/processor/sha_core/w[37] [12]),
	.F(\top/processor/sha_core/n3507_162 )
);
defparam \top/processor/sha_core/n3507_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_176 ),
	.I3(\top/processor/sha_core/n3507_161 ),
	.F(\top/processor/sha_core/n3879_124 )
);
defparam \top/processor/sha_core/n3879_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [12]),
	.I2(\top/processor/sha_core/w[39] [12]),
	.F(\top/processor/sha_core/n3879_125 )
);
defparam \top/processor/sha_core/n3879_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_127 ),
	.I3(\top/processor/sha_core/n3507_177 ),
	.F(\top/processor/sha_core/n3507_163 )
);
defparam \top/processor/sha_core/n3507_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [12]),
	.I2(\top/processor/sha_core/w[41] [12]),
	.F(\top/processor/sha_core/n3507_164 )
);
defparam \top/processor/sha_core/n3507_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [12]),
	.I2(\top/processor/sha_core/w[45] [12]),
	.F(\top/processor/sha_core/n3507_165 )
);
defparam \top/processor/sha_core/n3507_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_177 ),
	.I3(\top/processor/sha_core/n3507_164 ),
	.F(\top/processor/sha_core/n3879_126 )
);
defparam \top/processor/sha_core/n3879_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [12]),
	.I2(\top/processor/sha_core/w[47] [12]),
	.F(\top/processor/sha_core/n3879_127 )
);
defparam \top/processor/sha_core/n3879_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_129 ),
	.I3(\top/processor/sha_core/n3507_178 ),
	.F(\top/processor/sha_core/n3507_166 )
);
defparam \top/processor/sha_core/n3507_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [12]),
	.I2(\top/processor/sha_core/w[49] [12]),
	.F(\top/processor/sha_core/n3507_167 )
);
defparam \top/processor/sha_core/n3507_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [12]),
	.I2(\top/processor/sha_core/w[53] [12]),
	.F(\top/processor/sha_core/n3507_168 )
);
defparam \top/processor/sha_core/n3507_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_178 ),
	.I3(\top/processor/sha_core/n3507_167 ),
	.F(\top/processor/sha_core/n3879_128 )
);
defparam \top/processor/sha_core/n3879_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [12]),
	.I2(\top/processor/sha_core/w[55] [12]),
	.F(\top/processor/sha_core/n3879_129 )
);
defparam \top/processor/sha_core/n3879_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3507_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3879_131 ),
	.I3(\top/processor/sha_core/n3507_179 ),
	.F(\top/processor/sha_core/n3507_169 )
);
defparam \top/processor/sha_core/n3507_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3507_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [12]),
	.I2(\top/processor/sha_core/w[57] [12]),
	.F(\top/processor/sha_core/n3507_170 )
);
defparam \top/processor/sha_core/n3507_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [12]),
	.I2(\top/processor/sha_core/w[61] [12]),
	.F(\top/processor/sha_core/n3507_171 )
);
defparam \top/processor/sha_core/n3507_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3879_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3507_179 ),
	.I3(\top/processor/sha_core/n3507_170 ),
	.F(\top/processor/sha_core/n3879_130 )
);
defparam \top/processor/sha_core/n3879_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3879_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [12]),
	.I2(\top/processor/sha_core/w[63] [12]),
	.F(\top/processor/sha_core/n3879_131 )
);
defparam \top/processor/sha_core/n3879_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3489_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3861_131 ),
	.I3(\top/processor/sha_core/n3489_179 ),
	.F(\top/processor/sha_core/n3489_169 )
);
defparam \top/processor/sha_core/n3489_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3489_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [30]),
	.I2(\top/processor/sha_core/w[57] [30]),
	.F(\top/processor/sha_core/n3489_170 )
);
defparam \top/processor/sha_core/n3489_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [30]),
	.I2(\top/processor/sha_core/w[61] [30]),
	.F(\top/processor/sha_core/n3489_171 )
);
defparam \top/processor/sha_core/n3489_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3861_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3489_179 ),
	.I3(\top/processor/sha_core/n3489_170 ),
	.F(\top/processor/sha_core/n3861_130 )
);
defparam \top/processor/sha_core/n3861_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3861_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [30]),
	.I2(\top/processor/sha_core/w[63] [30]),
	.F(\top/processor/sha_core/n3861_131 )
);
defparam \top/processor/sha_core/n3861_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_117 ),
	.I3(\top/processor/sha_core/n3508_172 ),
	.F(\top/processor/sha_core/n3508_148 )
);
defparam \top/processor/sha_core/n3508_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [11]),
	.I2(\top/processor/sha_core/w[1] [11]),
	.F(\top/processor/sha_core/n3508_149 )
);
defparam \top/processor/sha_core/n3508_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [11]),
	.I2(\top/processor/sha_core/w[5] [11]),
	.F(\top/processor/sha_core/n3508_150 )
);
defparam \top/processor/sha_core/n3508_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_172 ),
	.I3(\top/processor/sha_core/n3508_149 ),
	.F(\top/processor/sha_core/n3880_116 )
);
defparam \top/processor/sha_core/n3880_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [11]),
	.I2(\top/processor/sha_core/w[7] [11]),
	.F(\top/processor/sha_core/n3880_117 )
);
defparam \top/processor/sha_core/n3880_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_119 ),
	.I3(\top/processor/sha_core/n3508_173 ),
	.F(\top/processor/sha_core/n3508_151 )
);
defparam \top/processor/sha_core/n3508_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [11]),
	.I2(\top/processor/sha_core/w[9] [11]),
	.F(\top/processor/sha_core/n3508_152 )
);
defparam \top/processor/sha_core/n3508_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [11]),
	.I2(\top/processor/sha_core/w[13] [11]),
	.F(\top/processor/sha_core/n3508_153 )
);
defparam \top/processor/sha_core/n3508_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_173 ),
	.I3(\top/processor/sha_core/n3508_152 ),
	.F(\top/processor/sha_core/n3880_118 )
);
defparam \top/processor/sha_core/n3880_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [11]),
	.I2(\top/processor/sha_core/w[15] [11]),
	.F(\top/processor/sha_core/n3880_119 )
);
defparam \top/processor/sha_core/n3880_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_121 ),
	.I3(\top/processor/sha_core/n3508_174 ),
	.F(\top/processor/sha_core/n3508_154 )
);
defparam \top/processor/sha_core/n3508_s141 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3508_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [11]),
	.I2(\top/processor/sha_core/w[17] [11]),
	.F(\top/processor/sha_core/n3508_155 )
);
defparam \top/processor/sha_core/n3508_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [11]),
	.I2(\top/processor/sha_core/w[21] [11]),
	.F(\top/processor/sha_core/n3508_156 )
);
defparam \top/processor/sha_core/n3508_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_174 ),
	.I3(\top/processor/sha_core/n3508_155 ),
	.F(\top/processor/sha_core/n3880_120 )
);
defparam \top/processor/sha_core/n3880_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [11]),
	.I2(\top/processor/sha_core/w[23] [11]),
	.F(\top/processor/sha_core/n3880_121 )
);
defparam \top/processor/sha_core/n3880_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_123 ),
	.I3(\top/processor/sha_core/n3508_175 ),
	.F(\top/processor/sha_core/n3508_157 )
);
defparam \top/processor/sha_core/n3508_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [11]),
	.I2(\top/processor/sha_core/w[25] [11]),
	.F(\top/processor/sha_core/n3508_158 )
);
defparam \top/processor/sha_core/n3508_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [11]),
	.I2(\top/processor/sha_core/w[29] [11]),
	.F(\top/processor/sha_core/n3508_159 )
);
defparam \top/processor/sha_core/n3508_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_175 ),
	.I3(\top/processor/sha_core/n3508_158 ),
	.F(\top/processor/sha_core/n3880_122 )
);
defparam \top/processor/sha_core/n3880_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [11]),
	.I2(\top/processor/sha_core/w[31] [11]),
	.F(\top/processor/sha_core/n3880_123 )
);
defparam \top/processor/sha_core/n3880_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_125 ),
	.I3(\top/processor/sha_core/n3508_176 ),
	.F(\top/processor/sha_core/n3508_160 )
);
defparam \top/processor/sha_core/n3508_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [11]),
	.I2(\top/processor/sha_core/w[33] [11]),
	.F(\top/processor/sha_core/n3508_161 )
);
defparam \top/processor/sha_core/n3508_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [11]),
	.I2(\top/processor/sha_core/w[37] [11]),
	.F(\top/processor/sha_core/n3508_162 )
);
defparam \top/processor/sha_core/n3508_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_176 ),
	.I3(\top/processor/sha_core/n3508_161 ),
	.F(\top/processor/sha_core/n3880_124 )
);
defparam \top/processor/sha_core/n3880_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [11]),
	.I2(\top/processor/sha_core/w[39] [11]),
	.F(\top/processor/sha_core/n3880_125 )
);
defparam \top/processor/sha_core/n3880_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_127 ),
	.I3(\top/processor/sha_core/n3508_177 ),
	.F(\top/processor/sha_core/n3508_163 )
);
defparam \top/processor/sha_core/n3508_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [11]),
	.I2(\top/processor/sha_core/w[41] [11]),
	.F(\top/processor/sha_core/n3508_164 )
);
defparam \top/processor/sha_core/n3508_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [11]),
	.I2(\top/processor/sha_core/w[45] [11]),
	.F(\top/processor/sha_core/n3508_165 )
);
defparam \top/processor/sha_core/n3508_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_177 ),
	.I3(\top/processor/sha_core/n3508_164 ),
	.F(\top/processor/sha_core/n3880_126 )
);
defparam \top/processor/sha_core/n3880_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [11]),
	.I2(\top/processor/sha_core/w[47] [11]),
	.F(\top/processor/sha_core/n3880_127 )
);
defparam \top/processor/sha_core/n3880_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_129 ),
	.I3(\top/processor/sha_core/n3508_178 ),
	.F(\top/processor/sha_core/n3508_166 )
);
defparam \top/processor/sha_core/n3508_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [11]),
	.I2(\top/processor/sha_core/w[49] [11]),
	.F(\top/processor/sha_core/n3508_167 )
);
defparam \top/processor/sha_core/n3508_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [11]),
	.I2(\top/processor/sha_core/w[53] [11]),
	.F(\top/processor/sha_core/n3508_168 )
);
defparam \top/processor/sha_core/n3508_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_178 ),
	.I3(\top/processor/sha_core/n3508_167 ),
	.F(\top/processor/sha_core/n3880_128 )
);
defparam \top/processor/sha_core/n3880_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3880_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [11]),
	.I2(\top/processor/sha_core/w[55] [11]),
	.F(\top/processor/sha_core/n3880_129 )
);
defparam \top/processor/sha_core/n3880_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3508_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3880_131 ),
	.I3(\top/processor/sha_core/n3508_179 ),
	.F(\top/processor/sha_core/n3508_169 )
);
defparam \top/processor/sha_core/n3508_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3508_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [11]),
	.I2(\top/processor/sha_core/w[57] [11]),
	.F(\top/processor/sha_core/n3508_170 )
);
defparam \top/processor/sha_core/n3508_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [11]),
	.I2(\top/processor/sha_core/w[61] [11]),
	.F(\top/processor/sha_core/n3508_171 )
);
defparam \top/processor/sha_core/n3508_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3880_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3508_179 ),
	.I3(\top/processor/sha_core/n3508_170 ),
	.F(\top/processor/sha_core/n3880_130 )
);
defparam \top/processor/sha_core/n3880_s117 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3880_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [11]),
	.I2(\top/processor/sha_core/w[63] [11]),
	.F(\top/processor/sha_core/n3880_131 )
);
defparam \top/processor/sha_core/n3880_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_117 ),
	.I3(\top/processor/sha_core/n3509_172 ),
	.F(\top/processor/sha_core/n3509_148 )
);
defparam \top/processor/sha_core/n3509_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [10]),
	.I2(\top/processor/sha_core/w[1] [10]),
	.F(\top/processor/sha_core/n3509_149 )
);
defparam \top/processor/sha_core/n3509_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [10]),
	.I2(\top/processor/sha_core/w[5] [10]),
	.F(\top/processor/sha_core/n3509_150 )
);
defparam \top/processor/sha_core/n3509_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_172 ),
	.I3(\top/processor/sha_core/n3509_149 ),
	.F(\top/processor/sha_core/n3881_116 )
);
defparam \top/processor/sha_core/n3881_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [10]),
	.I2(\top/processor/sha_core/w[7] [10]),
	.F(\top/processor/sha_core/n3881_117 )
);
defparam \top/processor/sha_core/n3881_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_119 ),
	.I3(\top/processor/sha_core/n3509_173 ),
	.F(\top/processor/sha_core/n3509_151 )
);
defparam \top/processor/sha_core/n3509_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [10]),
	.I2(\top/processor/sha_core/w[9] [10]),
	.F(\top/processor/sha_core/n3509_152 )
);
defparam \top/processor/sha_core/n3509_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [10]),
	.I2(\top/processor/sha_core/w[13] [10]),
	.F(\top/processor/sha_core/n3509_153 )
);
defparam \top/processor/sha_core/n3509_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_173 ),
	.I3(\top/processor/sha_core/n3509_152 ),
	.F(\top/processor/sha_core/n3881_118 )
);
defparam \top/processor/sha_core/n3881_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [10]),
	.I2(\top/processor/sha_core/w[15] [10]),
	.F(\top/processor/sha_core/n3881_119 )
);
defparam \top/processor/sha_core/n3881_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_117 ),
	.I3(\top/processor/sha_core/n3490_172 ),
	.F(\top/processor/sha_core/n3490_148 )
);
defparam \top/processor/sha_core/n3490_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [29]),
	.I2(\top/processor/sha_core/w[1] [29]),
	.F(\top/processor/sha_core/n3490_149 )
);
defparam \top/processor/sha_core/n3490_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [29]),
	.I2(\top/processor/sha_core/w[5] [29]),
	.F(\top/processor/sha_core/n3490_150 )
);
defparam \top/processor/sha_core/n3490_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_172 ),
	.I3(\top/processor/sha_core/n3490_149 ),
	.F(\top/processor/sha_core/n3862_116 )
);
defparam \top/processor/sha_core/n3862_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [29]),
	.I2(\top/processor/sha_core/w[7] [29]),
	.F(\top/processor/sha_core/n3862_117 )
);
defparam \top/processor/sha_core/n3862_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_121 ),
	.I3(\top/processor/sha_core/n3509_174 ),
	.F(\top/processor/sha_core/n3509_154 )
);
defparam \top/processor/sha_core/n3509_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [10]),
	.I2(\top/processor/sha_core/w[17] [10]),
	.F(\top/processor/sha_core/n3509_155 )
);
defparam \top/processor/sha_core/n3509_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [10]),
	.I2(\top/processor/sha_core/w[21] [10]),
	.F(\top/processor/sha_core/n3509_156 )
);
defparam \top/processor/sha_core/n3509_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_174 ),
	.I3(\top/processor/sha_core/n3509_155 ),
	.F(\top/processor/sha_core/n3881_120 )
);
defparam \top/processor/sha_core/n3881_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [10]),
	.I2(\top/processor/sha_core/w[23] [10]),
	.F(\top/processor/sha_core/n3881_121 )
);
defparam \top/processor/sha_core/n3881_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_123 ),
	.I3(\top/processor/sha_core/n3509_175 ),
	.F(\top/processor/sha_core/n3509_157 )
);
defparam \top/processor/sha_core/n3509_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [10]),
	.I2(\top/processor/sha_core/w[25] [10]),
	.F(\top/processor/sha_core/n3509_158 )
);
defparam \top/processor/sha_core/n3509_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [10]),
	.I2(\top/processor/sha_core/w[29] [10]),
	.F(\top/processor/sha_core/n3509_159 )
);
defparam \top/processor/sha_core/n3509_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_175 ),
	.I3(\top/processor/sha_core/n3509_158 ),
	.F(\top/processor/sha_core/n3881_122 )
);
defparam \top/processor/sha_core/n3881_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [10]),
	.I2(\top/processor/sha_core/w[31] [10]),
	.F(\top/processor/sha_core/n3881_123 )
);
defparam \top/processor/sha_core/n3881_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_125 ),
	.I3(\top/processor/sha_core/n3509_176 ),
	.F(\top/processor/sha_core/n3509_160 )
);
defparam \top/processor/sha_core/n3509_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [10]),
	.I2(\top/processor/sha_core/w[33] [10]),
	.F(\top/processor/sha_core/n3509_161 )
);
defparam \top/processor/sha_core/n3509_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [10]),
	.I2(\top/processor/sha_core/w[37] [10]),
	.F(\top/processor/sha_core/n3509_162 )
);
defparam \top/processor/sha_core/n3509_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_176 ),
	.I3(\top/processor/sha_core/n3509_161 ),
	.F(\top/processor/sha_core/n3881_124 )
);
defparam \top/processor/sha_core/n3881_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [10]),
	.I2(\top/processor/sha_core/w[39] [10]),
	.F(\top/processor/sha_core/n3881_125 )
);
defparam \top/processor/sha_core/n3881_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_127 ),
	.I3(\top/processor/sha_core/n3509_177 ),
	.F(\top/processor/sha_core/n3509_163 )
);
defparam \top/processor/sha_core/n3509_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [10]),
	.I2(\top/processor/sha_core/w[41] [10]),
	.F(\top/processor/sha_core/n3509_164 )
);
defparam \top/processor/sha_core/n3509_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [10]),
	.I2(\top/processor/sha_core/w[45] [10]),
	.F(\top/processor/sha_core/n3509_165 )
);
defparam \top/processor/sha_core/n3509_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_177 ),
	.I3(\top/processor/sha_core/n3509_164 ),
	.F(\top/processor/sha_core/n3881_126 )
);
defparam \top/processor/sha_core/n3881_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [10]),
	.I2(\top/processor/sha_core/w[47] [10]),
	.F(\top/processor/sha_core/n3881_127 )
);
defparam \top/processor/sha_core/n3881_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_129 ),
	.I3(\top/processor/sha_core/n3509_178 ),
	.F(\top/processor/sha_core/n3509_166 )
);
defparam \top/processor/sha_core/n3509_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [10]),
	.I2(\top/processor/sha_core/w[49] [10]),
	.F(\top/processor/sha_core/n3509_167 )
);
defparam \top/processor/sha_core/n3509_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [10]),
	.I2(\top/processor/sha_core/w[53] [10]),
	.F(\top/processor/sha_core/n3509_168 )
);
defparam \top/processor/sha_core/n3509_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_178 ),
	.I3(\top/processor/sha_core/n3509_167 ),
	.F(\top/processor/sha_core/n3881_128 )
);
defparam \top/processor/sha_core/n3881_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [10]),
	.I2(\top/processor/sha_core/w[55] [10]),
	.F(\top/processor/sha_core/n3881_129 )
);
defparam \top/processor/sha_core/n3881_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3509_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3881_131 ),
	.I3(\top/processor/sha_core/n3509_179 ),
	.F(\top/processor/sha_core/n3509_169 )
);
defparam \top/processor/sha_core/n3509_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3509_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [10]),
	.I2(\top/processor/sha_core/w[57] [10]),
	.F(\top/processor/sha_core/n3509_170 )
);
defparam \top/processor/sha_core/n3509_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [10]),
	.I2(\top/processor/sha_core/w[61] [10]),
	.F(\top/processor/sha_core/n3509_171 )
);
defparam \top/processor/sha_core/n3509_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3881_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3509_179 ),
	.I3(\top/processor/sha_core/n3509_170 ),
	.F(\top/processor/sha_core/n3881_130 )
);
defparam \top/processor/sha_core/n3881_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3881_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [10]),
	.I2(\top/processor/sha_core/w[63] [10]),
	.F(\top/processor/sha_core/n3881_131 )
);
defparam \top/processor/sha_core/n3881_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_117 ),
	.I3(\top/processor/sha_core/n3510_172 ),
	.F(\top/processor/sha_core/n3510_148 )
);
defparam \top/processor/sha_core/n3510_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [9]),
	.I2(\top/processor/sha_core/w[1] [9]),
	.F(\top/processor/sha_core/n3510_149 )
);
defparam \top/processor/sha_core/n3510_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [9]),
	.I2(\top/processor/sha_core/w[5] [9]),
	.F(\top/processor/sha_core/n3510_150 )
);
defparam \top/processor/sha_core/n3510_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_172 ),
	.I3(\top/processor/sha_core/n3510_149 ),
	.F(\top/processor/sha_core/n3882_116 )
);
defparam \top/processor/sha_core/n3882_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [9]),
	.I2(\top/processor/sha_core/w[7] [9]),
	.F(\top/processor/sha_core/n3882_117 )
);
defparam \top/processor/sha_core/n3882_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_119 ),
	.I3(\top/processor/sha_core/n3510_173 ),
	.F(\top/processor/sha_core/n3510_151 )
);
defparam \top/processor/sha_core/n3510_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [9]),
	.I2(\top/processor/sha_core/w[9] [9]),
	.F(\top/processor/sha_core/n3510_152 )
);
defparam \top/processor/sha_core/n3510_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [9]),
	.I2(\top/processor/sha_core/w[13] [9]),
	.F(\top/processor/sha_core/n3510_153 )
);
defparam \top/processor/sha_core/n3510_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_173 ),
	.I3(\top/processor/sha_core/n3510_152 ),
	.F(\top/processor/sha_core/n3882_118 )
);
defparam \top/processor/sha_core/n3882_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [9]),
	.I2(\top/processor/sha_core/w[15] [9]),
	.F(\top/processor/sha_core/n3882_119 )
);
defparam \top/processor/sha_core/n3882_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_121 ),
	.I3(\top/processor/sha_core/n3510_174 ),
	.F(\top/processor/sha_core/n3510_154 )
);
defparam \top/processor/sha_core/n3510_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [9]),
	.I2(\top/processor/sha_core/w[17] [9]),
	.F(\top/processor/sha_core/n3510_155 )
);
defparam \top/processor/sha_core/n3510_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [9]),
	.I2(\top/processor/sha_core/w[21] [9]),
	.F(\top/processor/sha_core/n3510_156 )
);
defparam \top/processor/sha_core/n3510_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_174 ),
	.I3(\top/processor/sha_core/n3510_155 ),
	.F(\top/processor/sha_core/n3882_120 )
);
defparam \top/processor/sha_core/n3882_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [9]),
	.I2(\top/processor/sha_core/w[23] [9]),
	.F(\top/processor/sha_core/n3882_121 )
);
defparam \top/processor/sha_core/n3882_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_123 ),
	.I3(\top/processor/sha_core/n3510_175 ),
	.F(\top/processor/sha_core/n3510_157 )
);
defparam \top/processor/sha_core/n3510_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [9]),
	.I2(\top/processor/sha_core/w[25] [9]),
	.F(\top/processor/sha_core/n3510_158 )
);
defparam \top/processor/sha_core/n3510_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [9]),
	.I2(\top/processor/sha_core/w[29] [9]),
	.F(\top/processor/sha_core/n3510_159 )
);
defparam \top/processor/sha_core/n3510_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_175 ),
	.I3(\top/processor/sha_core/n3510_158 ),
	.F(\top/processor/sha_core/n3882_122 )
);
defparam \top/processor/sha_core/n3882_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [9]),
	.I2(\top/processor/sha_core/w[31] [9]),
	.F(\top/processor/sha_core/n3882_123 )
);
defparam \top/processor/sha_core/n3882_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_119 ),
	.I3(\top/processor/sha_core/n3490_173 ),
	.F(\top/processor/sha_core/n3490_151 )
);
defparam \top/processor/sha_core/n3490_s138 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3490_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [29]),
	.I2(\top/processor/sha_core/w[9] [29]),
	.F(\top/processor/sha_core/n3490_152 )
);
defparam \top/processor/sha_core/n3490_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [29]),
	.I2(\top/processor/sha_core/w[13] [29]),
	.F(\top/processor/sha_core/n3490_153 )
);
defparam \top/processor/sha_core/n3490_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_173 ),
	.I3(\top/processor/sha_core/n3490_152 ),
	.F(\top/processor/sha_core/n3862_118 )
);
defparam \top/processor/sha_core/n3862_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [29]),
	.I2(\top/processor/sha_core/w[15] [29]),
	.F(\top/processor/sha_core/n3862_119 )
);
defparam \top/processor/sha_core/n3862_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_125 ),
	.I3(\top/processor/sha_core/n3510_176 ),
	.F(\top/processor/sha_core/n3510_160 )
);
defparam \top/processor/sha_core/n3510_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [9]),
	.I2(\top/processor/sha_core/w[33] [9]),
	.F(\top/processor/sha_core/n3510_161 )
);
defparam \top/processor/sha_core/n3510_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [9]),
	.I2(\top/processor/sha_core/w[37] [9]),
	.F(\top/processor/sha_core/n3510_162 )
);
defparam \top/processor/sha_core/n3510_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_176 ),
	.I3(\top/processor/sha_core/n3510_161 ),
	.F(\top/processor/sha_core/n3882_124 )
);
defparam \top/processor/sha_core/n3882_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [9]),
	.I2(\top/processor/sha_core/w[39] [9]),
	.F(\top/processor/sha_core/n3882_125 )
);
defparam \top/processor/sha_core/n3882_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_127 ),
	.I3(\top/processor/sha_core/n3510_177 ),
	.F(\top/processor/sha_core/n3510_163 )
);
defparam \top/processor/sha_core/n3510_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [9]),
	.I2(\top/processor/sha_core/w[41] [9]),
	.F(\top/processor/sha_core/n3510_164 )
);
defparam \top/processor/sha_core/n3510_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [9]),
	.I2(\top/processor/sha_core/w[45] [9]),
	.F(\top/processor/sha_core/n3510_165 )
);
defparam \top/processor/sha_core/n3510_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_177 ),
	.I3(\top/processor/sha_core/n3510_164 ),
	.F(\top/processor/sha_core/n3882_126 )
);
defparam \top/processor/sha_core/n3882_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [9]),
	.I2(\top/processor/sha_core/w[47] [9]),
	.F(\top/processor/sha_core/n3882_127 )
);
defparam \top/processor/sha_core/n3882_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_129 ),
	.I3(\top/processor/sha_core/n3510_178 ),
	.F(\top/processor/sha_core/n3510_166 )
);
defparam \top/processor/sha_core/n3510_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [9]),
	.I2(\top/processor/sha_core/w[49] [9]),
	.F(\top/processor/sha_core/n3510_167 )
);
defparam \top/processor/sha_core/n3510_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [9]),
	.I2(\top/processor/sha_core/w[53] [9]),
	.F(\top/processor/sha_core/n3510_168 )
);
defparam \top/processor/sha_core/n3510_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_178 ),
	.I3(\top/processor/sha_core/n3510_167 ),
	.F(\top/processor/sha_core/n3882_128 )
);
defparam \top/processor/sha_core/n3882_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [9]),
	.I2(\top/processor/sha_core/w[55] [9]),
	.F(\top/processor/sha_core/n3882_129 )
);
defparam \top/processor/sha_core/n3882_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3510_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3882_131 ),
	.I3(\top/processor/sha_core/n3510_179 ),
	.F(\top/processor/sha_core/n3510_169 )
);
defparam \top/processor/sha_core/n3510_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3510_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [9]),
	.I2(\top/processor/sha_core/w[57] [9]),
	.F(\top/processor/sha_core/n3510_170 )
);
defparam \top/processor/sha_core/n3510_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [9]),
	.I2(\top/processor/sha_core/w[61] [9]),
	.F(\top/processor/sha_core/n3510_171 )
);
defparam \top/processor/sha_core/n3510_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3882_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3510_179 ),
	.I3(\top/processor/sha_core/n3510_170 ),
	.F(\top/processor/sha_core/n3882_130 )
);
defparam \top/processor/sha_core/n3882_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3882_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [9]),
	.I2(\top/processor/sha_core/w[63] [9]),
	.F(\top/processor/sha_core/n3882_131 )
);
defparam \top/processor/sha_core/n3882_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_117 ),
	.I3(\top/processor/sha_core/n3511_172 ),
	.F(\top/processor/sha_core/n3511_148 )
);
defparam \top/processor/sha_core/n3511_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [8]),
	.I2(\top/processor/sha_core/w[1] [8]),
	.F(\top/processor/sha_core/n3511_149 )
);
defparam \top/processor/sha_core/n3511_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [8]),
	.I2(\top/processor/sha_core/w[5] [8]),
	.F(\top/processor/sha_core/n3511_150 )
);
defparam \top/processor/sha_core/n3511_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_172 ),
	.I3(\top/processor/sha_core/n3511_149 ),
	.F(\top/processor/sha_core/n3883_116 )
);
defparam \top/processor/sha_core/n3883_s103 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3883_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [8]),
	.I2(\top/processor/sha_core/w[7] [8]),
	.F(\top/processor/sha_core/n3883_117 )
);
defparam \top/processor/sha_core/n3883_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_119 ),
	.I3(\top/processor/sha_core/n3511_173 ),
	.F(\top/processor/sha_core/n3511_151 )
);
defparam \top/processor/sha_core/n3511_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [8]),
	.I2(\top/processor/sha_core/w[9] [8]),
	.F(\top/processor/sha_core/n3511_152 )
);
defparam \top/processor/sha_core/n3511_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [8]),
	.I2(\top/processor/sha_core/w[13] [8]),
	.F(\top/processor/sha_core/n3511_153 )
);
defparam \top/processor/sha_core/n3511_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_173 ),
	.I3(\top/processor/sha_core/n3511_152 ),
	.F(\top/processor/sha_core/n3883_118 )
);
defparam \top/processor/sha_core/n3883_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [8]),
	.I2(\top/processor/sha_core/w[15] [8]),
	.F(\top/processor/sha_core/n3883_119 )
);
defparam \top/processor/sha_core/n3883_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_121 ),
	.I3(\top/processor/sha_core/n3511_174 ),
	.F(\top/processor/sha_core/n3511_154 )
);
defparam \top/processor/sha_core/n3511_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [8]),
	.I2(\top/processor/sha_core/w[17] [8]),
	.F(\top/processor/sha_core/n3511_155 )
);
defparam \top/processor/sha_core/n3511_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [8]),
	.I2(\top/processor/sha_core/w[21] [8]),
	.F(\top/processor/sha_core/n3511_156 )
);
defparam \top/processor/sha_core/n3511_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_174 ),
	.I3(\top/processor/sha_core/n3511_155 ),
	.F(\top/processor/sha_core/n3883_120 )
);
defparam \top/processor/sha_core/n3883_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [8]),
	.I2(\top/processor/sha_core/w[23] [8]),
	.F(\top/processor/sha_core/n3883_121 )
);
defparam \top/processor/sha_core/n3883_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_123 ),
	.I3(\top/processor/sha_core/n3511_175 ),
	.F(\top/processor/sha_core/n3511_157 )
);
defparam \top/processor/sha_core/n3511_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [8]),
	.I2(\top/processor/sha_core/w[25] [8]),
	.F(\top/processor/sha_core/n3511_158 )
);
defparam \top/processor/sha_core/n3511_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [8]),
	.I2(\top/processor/sha_core/w[29] [8]),
	.F(\top/processor/sha_core/n3511_159 )
);
defparam \top/processor/sha_core/n3511_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_175 ),
	.I3(\top/processor/sha_core/n3511_158 ),
	.F(\top/processor/sha_core/n3883_122 )
);
defparam \top/processor/sha_core/n3883_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [8]),
	.I2(\top/processor/sha_core/w[31] [8]),
	.F(\top/processor/sha_core/n3883_123 )
);
defparam \top/processor/sha_core/n3883_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_125 ),
	.I3(\top/processor/sha_core/n3511_176 ),
	.F(\top/processor/sha_core/n3511_160 )
);
defparam \top/processor/sha_core/n3511_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [8]),
	.I2(\top/processor/sha_core/w[33] [8]),
	.F(\top/processor/sha_core/n3511_161 )
);
defparam \top/processor/sha_core/n3511_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [8]),
	.I2(\top/processor/sha_core/w[37] [8]),
	.F(\top/processor/sha_core/n3511_162 )
);
defparam \top/processor/sha_core/n3511_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_176 ),
	.I3(\top/processor/sha_core/n3511_161 ),
	.F(\top/processor/sha_core/n3883_124 )
);
defparam \top/processor/sha_core/n3883_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [8]),
	.I2(\top/processor/sha_core/w[39] [8]),
	.F(\top/processor/sha_core/n3883_125 )
);
defparam \top/processor/sha_core/n3883_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_127 ),
	.I3(\top/processor/sha_core/n3511_177 ),
	.F(\top/processor/sha_core/n3511_163 )
);
defparam \top/processor/sha_core/n3511_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [8]),
	.I2(\top/processor/sha_core/w[41] [8]),
	.F(\top/processor/sha_core/n3511_164 )
);
defparam \top/processor/sha_core/n3511_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [8]),
	.I2(\top/processor/sha_core/w[45] [8]),
	.F(\top/processor/sha_core/n3511_165 )
);
defparam \top/processor/sha_core/n3511_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_177 ),
	.I3(\top/processor/sha_core/n3511_164 ),
	.F(\top/processor/sha_core/n3883_126 )
);
defparam \top/processor/sha_core/n3883_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [8]),
	.I2(\top/processor/sha_core/w[47] [8]),
	.F(\top/processor/sha_core/n3883_127 )
);
defparam \top/processor/sha_core/n3883_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_121 ),
	.I3(\top/processor/sha_core/n3490_174 ),
	.F(\top/processor/sha_core/n3490_154 )
);
defparam \top/processor/sha_core/n3490_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [29]),
	.I2(\top/processor/sha_core/w[17] [29]),
	.F(\top/processor/sha_core/n3490_155 )
);
defparam \top/processor/sha_core/n3490_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [29]),
	.I2(\top/processor/sha_core/w[21] [29]),
	.F(\top/processor/sha_core/n3490_156 )
);
defparam \top/processor/sha_core/n3490_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_174 ),
	.I3(\top/processor/sha_core/n3490_155 ),
	.F(\top/processor/sha_core/n3862_120 )
);
defparam \top/processor/sha_core/n3862_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [29]),
	.I2(\top/processor/sha_core/w[23] [29]),
	.F(\top/processor/sha_core/n3862_121 )
);
defparam \top/processor/sha_core/n3862_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_129 ),
	.I3(\top/processor/sha_core/n3511_178 ),
	.F(\top/processor/sha_core/n3511_166 )
);
defparam \top/processor/sha_core/n3511_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [8]),
	.I2(\top/processor/sha_core/w[49] [8]),
	.F(\top/processor/sha_core/n3511_167 )
);
defparam \top/processor/sha_core/n3511_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [8]),
	.I2(\top/processor/sha_core/w[53] [8]),
	.F(\top/processor/sha_core/n3511_168 )
);
defparam \top/processor/sha_core/n3511_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_178 ),
	.I3(\top/processor/sha_core/n3511_167 ),
	.F(\top/processor/sha_core/n3883_128 )
);
defparam \top/processor/sha_core/n3883_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [8]),
	.I2(\top/processor/sha_core/w[55] [8]),
	.F(\top/processor/sha_core/n3883_129 )
);
defparam \top/processor/sha_core/n3883_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3511_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3883_131 ),
	.I3(\top/processor/sha_core/n3511_179 ),
	.F(\top/processor/sha_core/n3511_169 )
);
defparam \top/processor/sha_core/n3511_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3511_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [8]),
	.I2(\top/processor/sha_core/w[57] [8]),
	.F(\top/processor/sha_core/n3511_170 )
);
defparam \top/processor/sha_core/n3511_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [8]),
	.I2(\top/processor/sha_core/w[61] [8]),
	.F(\top/processor/sha_core/n3511_171 )
);
defparam \top/processor/sha_core/n3511_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3883_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3511_179 ),
	.I3(\top/processor/sha_core/n3511_170 ),
	.F(\top/processor/sha_core/n3883_130 )
);
defparam \top/processor/sha_core/n3883_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3883_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [8]),
	.I2(\top/processor/sha_core/w[63] [8]),
	.F(\top/processor/sha_core/n3883_131 )
);
defparam \top/processor/sha_core/n3883_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_117 ),
	.I3(\top/processor/sha_core/n3512_172 ),
	.F(\top/processor/sha_core/n3512_148 )
);
defparam \top/processor/sha_core/n3512_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [7]),
	.I2(\top/processor/sha_core/w[1] [7]),
	.F(\top/processor/sha_core/n3512_149 )
);
defparam \top/processor/sha_core/n3512_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [7]),
	.I2(\top/processor/sha_core/w[5] [7]),
	.F(\top/processor/sha_core/n3512_150 )
);
defparam \top/processor/sha_core/n3512_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_172 ),
	.I3(\top/processor/sha_core/n3512_149 ),
	.F(\top/processor/sha_core/n3884_116 )
);
defparam \top/processor/sha_core/n3884_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [7]),
	.I2(\top/processor/sha_core/w[7] [7]),
	.F(\top/processor/sha_core/n3884_117 )
);
defparam \top/processor/sha_core/n3884_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_119 ),
	.I3(\top/processor/sha_core/n3512_173 ),
	.F(\top/processor/sha_core/n3512_151 )
);
defparam \top/processor/sha_core/n3512_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [7]),
	.I2(\top/processor/sha_core/w[9] [7]),
	.F(\top/processor/sha_core/n3512_152 )
);
defparam \top/processor/sha_core/n3512_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [7]),
	.I2(\top/processor/sha_core/w[13] [7]),
	.F(\top/processor/sha_core/n3512_153 )
);
defparam \top/processor/sha_core/n3512_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_173 ),
	.I3(\top/processor/sha_core/n3512_152 ),
	.F(\top/processor/sha_core/n3884_118 )
);
defparam \top/processor/sha_core/n3884_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [7]),
	.I2(\top/processor/sha_core/w[15] [7]),
	.F(\top/processor/sha_core/n3884_119 )
);
defparam \top/processor/sha_core/n3884_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_121 ),
	.I3(\top/processor/sha_core/n3512_174 ),
	.F(\top/processor/sha_core/n3512_154 )
);
defparam \top/processor/sha_core/n3512_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [7]),
	.I2(\top/processor/sha_core/w[17] [7]),
	.F(\top/processor/sha_core/n3512_155 )
);
defparam \top/processor/sha_core/n3512_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [7]),
	.I2(\top/processor/sha_core/w[21] [7]),
	.F(\top/processor/sha_core/n3512_156 )
);
defparam \top/processor/sha_core/n3512_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_174 ),
	.I3(\top/processor/sha_core/n3512_155 ),
	.F(\top/processor/sha_core/n3884_120 )
);
defparam \top/processor/sha_core/n3884_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [7]),
	.I2(\top/processor/sha_core/w[23] [7]),
	.F(\top/processor/sha_core/n3884_121 )
);
defparam \top/processor/sha_core/n3884_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_123 ),
	.I3(\top/processor/sha_core/n3512_175 ),
	.F(\top/processor/sha_core/n3512_157 )
);
defparam \top/processor/sha_core/n3512_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [7]),
	.I2(\top/processor/sha_core/w[25] [7]),
	.F(\top/processor/sha_core/n3512_158 )
);
defparam \top/processor/sha_core/n3512_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [7]),
	.I2(\top/processor/sha_core/w[29] [7]),
	.F(\top/processor/sha_core/n3512_159 )
);
defparam \top/processor/sha_core/n3512_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_175 ),
	.I3(\top/processor/sha_core/n3512_158 ),
	.F(\top/processor/sha_core/n3884_122 )
);
defparam \top/processor/sha_core/n3884_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [7]),
	.I2(\top/processor/sha_core/w[31] [7]),
	.F(\top/processor/sha_core/n3884_123 )
);
defparam \top/processor/sha_core/n3884_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_125 ),
	.I3(\top/processor/sha_core/n3512_176 ),
	.F(\top/processor/sha_core/n3512_160 )
);
defparam \top/processor/sha_core/n3512_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [7]),
	.I2(\top/processor/sha_core/w[33] [7]),
	.F(\top/processor/sha_core/n3512_161 )
);
defparam \top/processor/sha_core/n3512_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [7]),
	.I2(\top/processor/sha_core/w[37] [7]),
	.F(\top/processor/sha_core/n3512_162 )
);
defparam \top/processor/sha_core/n3512_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_176 ),
	.I3(\top/processor/sha_core/n3512_161 ),
	.F(\top/processor/sha_core/n3884_124 )
);
defparam \top/processor/sha_core/n3884_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [7]),
	.I2(\top/processor/sha_core/w[39] [7]),
	.F(\top/processor/sha_core/n3884_125 )
);
defparam \top/processor/sha_core/n3884_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_127 ),
	.I3(\top/processor/sha_core/n3512_177 ),
	.F(\top/processor/sha_core/n3512_163 )
);
defparam \top/processor/sha_core/n3512_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [7]),
	.I2(\top/processor/sha_core/w[41] [7]),
	.F(\top/processor/sha_core/n3512_164 )
);
defparam \top/processor/sha_core/n3512_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [7]),
	.I2(\top/processor/sha_core/w[45] [7]),
	.F(\top/processor/sha_core/n3512_165 )
);
defparam \top/processor/sha_core/n3512_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_177 ),
	.I3(\top/processor/sha_core/n3512_164 ),
	.F(\top/processor/sha_core/n3884_126 )
);
defparam \top/processor/sha_core/n3884_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [7]),
	.I2(\top/processor/sha_core/w[47] [7]),
	.F(\top/processor/sha_core/n3884_127 )
);
defparam \top/processor/sha_core/n3884_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_129 ),
	.I3(\top/processor/sha_core/n3512_178 ),
	.F(\top/processor/sha_core/n3512_166 )
);
defparam \top/processor/sha_core/n3512_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [7]),
	.I2(\top/processor/sha_core/w[49] [7]),
	.F(\top/processor/sha_core/n3512_167 )
);
defparam \top/processor/sha_core/n3512_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [7]),
	.I2(\top/processor/sha_core/w[53] [7]),
	.F(\top/processor/sha_core/n3512_168 )
);
defparam \top/processor/sha_core/n3512_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_178 ),
	.I3(\top/processor/sha_core/n3512_167 ),
	.F(\top/processor/sha_core/n3884_128 )
);
defparam \top/processor/sha_core/n3884_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [7]),
	.I2(\top/processor/sha_core/w[55] [7]),
	.F(\top/processor/sha_core/n3884_129 )
);
defparam \top/processor/sha_core/n3884_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3512_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3884_131 ),
	.I3(\top/processor/sha_core/n3512_179 ),
	.F(\top/processor/sha_core/n3512_169 )
);
defparam \top/processor/sha_core/n3512_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3512_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [7]),
	.I2(\top/processor/sha_core/w[57] [7]),
	.F(\top/processor/sha_core/n3512_170 )
);
defparam \top/processor/sha_core/n3512_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [7]),
	.I2(\top/processor/sha_core/w[61] [7]),
	.F(\top/processor/sha_core/n3512_171 )
);
defparam \top/processor/sha_core/n3512_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3884_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3512_179 ),
	.I3(\top/processor/sha_core/n3512_170 ),
	.F(\top/processor/sha_core/n3884_130 )
);
defparam \top/processor/sha_core/n3884_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3884_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [7]),
	.I2(\top/processor/sha_core/w[63] [7]),
	.F(\top/processor/sha_core/n3884_131 )
);
defparam \top/processor/sha_core/n3884_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_123 ),
	.I3(\top/processor/sha_core/n3490_175 ),
	.F(\top/processor/sha_core/n3490_157 )
);
defparam \top/processor/sha_core/n3490_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [29]),
	.I2(\top/processor/sha_core/w[25] [29]),
	.F(\top/processor/sha_core/n3490_158 )
);
defparam \top/processor/sha_core/n3490_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [29]),
	.I2(\top/processor/sha_core/w[29] [29]),
	.F(\top/processor/sha_core/n3490_159 )
);
defparam \top/processor/sha_core/n3490_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_175 ),
	.I3(\top/processor/sha_core/n3490_158 ),
	.F(\top/processor/sha_core/n3862_122 )
);
defparam \top/processor/sha_core/n3862_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [29]),
	.I2(\top/processor/sha_core/w[31] [29]),
	.F(\top/processor/sha_core/n3862_123 )
);
defparam \top/processor/sha_core/n3862_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_125 ),
	.I3(\top/processor/sha_core/n3488_176 ),
	.F(\top/processor/sha_core/n3488_160 )
);
defparam \top/processor/sha_core/n3488_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [31]),
	.I2(\top/processor/sha_core/w[9] [31]),
	.F(\top/processor/sha_core/n3488_161 )
);
defparam \top/processor/sha_core/n3488_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [31]),
	.I2(\top/processor/sha_core/w[13] [31]),
	.F(\top/processor/sha_core/n3488_162 )
);
defparam \top/processor/sha_core/n3488_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_176 ),
	.I3(\top/processor/sha_core/n3488_161 ),
	.F(\top/processor/sha_core/n3860_124 )
);
defparam \top/processor/sha_core/n3860_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [31]),
	.I2(\top/processor/sha_core/w[15] [31]),
	.F(\top/processor/sha_core/n3860_125 )
);
defparam \top/processor/sha_core/n3860_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_117 ),
	.I3(\top/processor/sha_core/n3513_172 ),
	.F(\top/processor/sha_core/n3513_148 )
);
defparam \top/processor/sha_core/n3513_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [6]),
	.I2(\top/processor/sha_core/w[1] [6]),
	.F(\top/processor/sha_core/n3513_149 )
);
defparam \top/processor/sha_core/n3513_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [6]),
	.I2(\top/processor/sha_core/w[5] [6]),
	.F(\top/processor/sha_core/n3513_150 )
);
defparam \top/processor/sha_core/n3513_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_172 ),
	.I3(\top/processor/sha_core/n3513_149 ),
	.F(\top/processor/sha_core/n3885_116 )
);
defparam \top/processor/sha_core/n3885_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [6]),
	.I2(\top/processor/sha_core/w[7] [6]),
	.F(\top/processor/sha_core/n3885_117 )
);
defparam \top/processor/sha_core/n3885_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_119 ),
	.I3(\top/processor/sha_core/n3513_173 ),
	.F(\top/processor/sha_core/n3513_151 )
);
defparam \top/processor/sha_core/n3513_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [6]),
	.I2(\top/processor/sha_core/w[9] [6]),
	.F(\top/processor/sha_core/n3513_152 )
);
defparam \top/processor/sha_core/n3513_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [6]),
	.I2(\top/processor/sha_core/w[13] [6]),
	.F(\top/processor/sha_core/n3513_153 )
);
defparam \top/processor/sha_core/n3513_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_173 ),
	.I3(\top/processor/sha_core/n3513_152 ),
	.F(\top/processor/sha_core/n3885_118 )
);
defparam \top/processor/sha_core/n3885_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [6]),
	.I2(\top/processor/sha_core/w[15] [6]),
	.F(\top/processor/sha_core/n3885_119 )
);
defparam \top/processor/sha_core/n3885_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_121 ),
	.I3(\top/processor/sha_core/n3513_174 ),
	.F(\top/processor/sha_core/n3513_154 )
);
defparam \top/processor/sha_core/n3513_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [6]),
	.I2(\top/processor/sha_core/w[17] [6]),
	.F(\top/processor/sha_core/n3513_155 )
);
defparam \top/processor/sha_core/n3513_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [6]),
	.I2(\top/processor/sha_core/w[21] [6]),
	.F(\top/processor/sha_core/n3513_156 )
);
defparam \top/processor/sha_core/n3513_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_174 ),
	.I3(\top/processor/sha_core/n3513_155 ),
	.F(\top/processor/sha_core/n3885_120 )
);
defparam \top/processor/sha_core/n3885_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [6]),
	.I2(\top/processor/sha_core/w[23] [6]),
	.F(\top/processor/sha_core/n3885_121 )
);
defparam \top/processor/sha_core/n3885_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_123 ),
	.I3(\top/processor/sha_core/n3513_175 ),
	.F(\top/processor/sha_core/n3513_157 )
);
defparam \top/processor/sha_core/n3513_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [6]),
	.I2(\top/processor/sha_core/w[25] [6]),
	.F(\top/processor/sha_core/n3513_158 )
);
defparam \top/processor/sha_core/n3513_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [6]),
	.I2(\top/processor/sha_core/w[29] [6]),
	.F(\top/processor/sha_core/n3513_159 )
);
defparam \top/processor/sha_core/n3513_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_175 ),
	.I3(\top/processor/sha_core/n3513_158 ),
	.F(\top/processor/sha_core/n3885_122 )
);
defparam \top/processor/sha_core/n3885_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [6]),
	.I2(\top/processor/sha_core/w[31] [6]),
	.F(\top/processor/sha_core/n3885_123 )
);
defparam \top/processor/sha_core/n3885_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_125 ),
	.I3(\top/processor/sha_core/n3513_176 ),
	.F(\top/processor/sha_core/n3513_160 )
);
defparam \top/processor/sha_core/n3513_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [6]),
	.I2(\top/processor/sha_core/w[33] [6]),
	.F(\top/processor/sha_core/n3513_161 )
);
defparam \top/processor/sha_core/n3513_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [6]),
	.I2(\top/processor/sha_core/w[37] [6]),
	.F(\top/processor/sha_core/n3513_162 )
);
defparam \top/processor/sha_core/n3513_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_176 ),
	.I3(\top/processor/sha_core/n3513_161 ),
	.F(\top/processor/sha_core/n3885_124 )
);
defparam \top/processor/sha_core/n3885_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [6]),
	.I2(\top/processor/sha_core/w[39] [6]),
	.F(\top/processor/sha_core/n3885_125 )
);
defparam \top/processor/sha_core/n3885_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_127 ),
	.I3(\top/processor/sha_core/n3513_177 ),
	.F(\top/processor/sha_core/n3513_163 )
);
defparam \top/processor/sha_core/n3513_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [6]),
	.I2(\top/processor/sha_core/w[41] [6]),
	.F(\top/processor/sha_core/n3513_164 )
);
defparam \top/processor/sha_core/n3513_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [6]),
	.I2(\top/processor/sha_core/w[45] [6]),
	.F(\top/processor/sha_core/n3513_165 )
);
defparam \top/processor/sha_core/n3513_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_177 ),
	.I3(\top/processor/sha_core/n3513_164 ),
	.F(\top/processor/sha_core/n3885_126 )
);
defparam \top/processor/sha_core/n3885_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [6]),
	.I2(\top/processor/sha_core/w[47] [6]),
	.F(\top/processor/sha_core/n3885_127 )
);
defparam \top/processor/sha_core/n3885_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_129 ),
	.I3(\top/processor/sha_core/n3513_178 ),
	.F(\top/processor/sha_core/n3513_166 )
);
defparam \top/processor/sha_core/n3513_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [6]),
	.I2(\top/processor/sha_core/w[49] [6]),
	.F(\top/processor/sha_core/n3513_167 )
);
defparam \top/processor/sha_core/n3513_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [6]),
	.I2(\top/processor/sha_core/w[53] [6]),
	.F(\top/processor/sha_core/n3513_168 )
);
defparam \top/processor/sha_core/n3513_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_178 ),
	.I3(\top/processor/sha_core/n3513_167 ),
	.F(\top/processor/sha_core/n3885_128 )
);
defparam \top/processor/sha_core/n3885_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [6]),
	.I2(\top/processor/sha_core/w[55] [6]),
	.F(\top/processor/sha_core/n3885_129 )
);
defparam \top/processor/sha_core/n3885_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3513_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3885_131 ),
	.I3(\top/processor/sha_core/n3513_179 ),
	.F(\top/processor/sha_core/n3513_169 )
);
defparam \top/processor/sha_core/n3513_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3513_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [6]),
	.I2(\top/processor/sha_core/w[57] [6]),
	.F(\top/processor/sha_core/n3513_170 )
);
defparam \top/processor/sha_core/n3513_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [6]),
	.I2(\top/processor/sha_core/w[61] [6]),
	.F(\top/processor/sha_core/n3513_171 )
);
defparam \top/processor/sha_core/n3513_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3885_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3513_179 ),
	.I3(\top/processor/sha_core/n3513_170 ),
	.F(\top/processor/sha_core/n3885_130 )
);
defparam \top/processor/sha_core/n3885_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3885_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [6]),
	.I2(\top/processor/sha_core/w[63] [6]),
	.F(\top/processor/sha_core/n3885_131 )
);
defparam \top/processor/sha_core/n3885_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_117 ),
	.I3(\top/processor/sha_core/n3514_172 ),
	.F(\top/processor/sha_core/n3514_148 )
);
defparam \top/processor/sha_core/n3514_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [5]),
	.I2(\top/processor/sha_core/w[1] [5]),
	.F(\top/processor/sha_core/n3514_149 )
);
defparam \top/processor/sha_core/n3514_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [5]),
	.I2(\top/processor/sha_core/w[5] [5]),
	.F(\top/processor/sha_core/n3514_150 )
);
defparam \top/processor/sha_core/n3514_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_172 ),
	.I3(\top/processor/sha_core/n3514_149 ),
	.F(\top/processor/sha_core/n3886_116 )
);
defparam \top/processor/sha_core/n3886_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [5]),
	.I2(\top/processor/sha_core/w[7] [5]),
	.F(\top/processor/sha_core/n3886_117 )
);
defparam \top/processor/sha_core/n3886_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_119 ),
	.I3(\top/processor/sha_core/n3514_173 ),
	.F(\top/processor/sha_core/n3514_151 )
);
defparam \top/processor/sha_core/n3514_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [5]),
	.I2(\top/processor/sha_core/w[9] [5]),
	.F(\top/processor/sha_core/n3514_152 )
);
defparam \top/processor/sha_core/n3514_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [5]),
	.I2(\top/processor/sha_core/w[13] [5]),
	.F(\top/processor/sha_core/n3514_153 )
);
defparam \top/processor/sha_core/n3514_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_173 ),
	.I3(\top/processor/sha_core/n3514_152 ),
	.F(\top/processor/sha_core/n3886_118 )
);
defparam \top/processor/sha_core/n3886_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [5]),
	.I2(\top/processor/sha_core/w[15] [5]),
	.F(\top/processor/sha_core/n3886_119 )
);
defparam \top/processor/sha_core/n3886_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_125 ),
	.I3(\top/processor/sha_core/n3490_176 ),
	.F(\top/processor/sha_core/n3490_160 )
);
defparam \top/processor/sha_core/n3490_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [29]),
	.I2(\top/processor/sha_core/w[33] [29]),
	.F(\top/processor/sha_core/n3490_161 )
);
defparam \top/processor/sha_core/n3490_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [29]),
	.I2(\top/processor/sha_core/w[37] [29]),
	.F(\top/processor/sha_core/n3490_162 )
);
defparam \top/processor/sha_core/n3490_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_176 ),
	.I3(\top/processor/sha_core/n3490_161 ),
	.F(\top/processor/sha_core/n3862_124 )
);
defparam \top/processor/sha_core/n3862_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [29]),
	.I2(\top/processor/sha_core/w[39] [29]),
	.F(\top/processor/sha_core/n3862_125 )
);
defparam \top/processor/sha_core/n3862_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_121 ),
	.I3(\top/processor/sha_core/n3514_174 ),
	.F(\top/processor/sha_core/n3514_154 )
);
defparam \top/processor/sha_core/n3514_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [5]),
	.I2(\top/processor/sha_core/w[17] [5]),
	.F(\top/processor/sha_core/n3514_155 )
);
defparam \top/processor/sha_core/n3514_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [5]),
	.I2(\top/processor/sha_core/w[21] [5]),
	.F(\top/processor/sha_core/n3514_156 )
);
defparam \top/processor/sha_core/n3514_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_174 ),
	.I3(\top/processor/sha_core/n3514_155 ),
	.F(\top/processor/sha_core/n3886_120 )
);
defparam \top/processor/sha_core/n3886_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [5]),
	.I2(\top/processor/sha_core/w[23] [5]),
	.F(\top/processor/sha_core/n3886_121 )
);
defparam \top/processor/sha_core/n3886_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_123 ),
	.I3(\top/processor/sha_core/n3514_175 ),
	.F(\top/processor/sha_core/n3514_157 )
);
defparam \top/processor/sha_core/n3514_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [5]),
	.I2(\top/processor/sha_core/w[25] [5]),
	.F(\top/processor/sha_core/n3514_158 )
);
defparam \top/processor/sha_core/n3514_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [5]),
	.I2(\top/processor/sha_core/w[29] [5]),
	.F(\top/processor/sha_core/n3514_159 )
);
defparam \top/processor/sha_core/n3514_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_175 ),
	.I3(\top/processor/sha_core/n3514_158 ),
	.F(\top/processor/sha_core/n3886_122 )
);
defparam \top/processor/sha_core/n3886_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [5]),
	.I2(\top/processor/sha_core/w[31] [5]),
	.F(\top/processor/sha_core/n3886_123 )
);
defparam \top/processor/sha_core/n3886_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_125 ),
	.I3(\top/processor/sha_core/n3514_176 ),
	.F(\top/processor/sha_core/n3514_160 )
);
defparam \top/processor/sha_core/n3514_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [5]),
	.I2(\top/processor/sha_core/w[33] [5]),
	.F(\top/processor/sha_core/n3514_161 )
);
defparam \top/processor/sha_core/n3514_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [5]),
	.I2(\top/processor/sha_core/w[37] [5]),
	.F(\top/processor/sha_core/n3514_162 )
);
defparam \top/processor/sha_core/n3514_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_176 ),
	.I3(\top/processor/sha_core/n3514_161 ),
	.F(\top/processor/sha_core/n3886_124 )
);
defparam \top/processor/sha_core/n3886_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [5]),
	.I2(\top/processor/sha_core/w[39] [5]),
	.F(\top/processor/sha_core/n3886_125 )
);
defparam \top/processor/sha_core/n3886_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_127 ),
	.I3(\top/processor/sha_core/n3514_177 ),
	.F(\top/processor/sha_core/n3514_163 )
);
defparam \top/processor/sha_core/n3514_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [5]),
	.I2(\top/processor/sha_core/w[41] [5]),
	.F(\top/processor/sha_core/n3514_164 )
);
defparam \top/processor/sha_core/n3514_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [5]),
	.I2(\top/processor/sha_core/w[45] [5]),
	.F(\top/processor/sha_core/n3514_165 )
);
defparam \top/processor/sha_core/n3514_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_177 ),
	.I3(\top/processor/sha_core/n3514_164 ),
	.F(\top/processor/sha_core/n3886_126 )
);
defparam \top/processor/sha_core/n3886_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [5]),
	.I2(\top/processor/sha_core/w[47] [5]),
	.F(\top/processor/sha_core/n3886_127 )
);
defparam \top/processor/sha_core/n3886_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_129 ),
	.I3(\top/processor/sha_core/n3514_178 ),
	.F(\top/processor/sha_core/n3514_166 )
);
defparam \top/processor/sha_core/n3514_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [5]),
	.I2(\top/processor/sha_core/w[49] [5]),
	.F(\top/processor/sha_core/n3514_167 )
);
defparam \top/processor/sha_core/n3514_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [5]),
	.I2(\top/processor/sha_core/w[53] [5]),
	.F(\top/processor/sha_core/n3514_168 )
);
defparam \top/processor/sha_core/n3514_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_178 ),
	.I3(\top/processor/sha_core/n3514_167 ),
	.F(\top/processor/sha_core/n3886_128 )
);
defparam \top/processor/sha_core/n3886_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [5]),
	.I2(\top/processor/sha_core/w[55] [5]),
	.F(\top/processor/sha_core/n3886_129 )
);
defparam \top/processor/sha_core/n3886_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3514_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3886_131 ),
	.I3(\top/processor/sha_core/n3514_179 ),
	.F(\top/processor/sha_core/n3514_169 )
);
defparam \top/processor/sha_core/n3514_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3514_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [5]),
	.I2(\top/processor/sha_core/w[57] [5]),
	.F(\top/processor/sha_core/n3514_170 )
);
defparam \top/processor/sha_core/n3514_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [5]),
	.I2(\top/processor/sha_core/w[61] [5]),
	.F(\top/processor/sha_core/n3514_171 )
);
defparam \top/processor/sha_core/n3514_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3886_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3514_179 ),
	.I3(\top/processor/sha_core/n3514_170 ),
	.F(\top/processor/sha_core/n3886_130 )
);
defparam \top/processor/sha_core/n3886_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3886_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [5]),
	.I2(\top/processor/sha_core/w[63] [5]),
	.F(\top/processor/sha_core/n3886_131 )
);
defparam \top/processor/sha_core/n3886_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_117 ),
	.I3(\top/processor/sha_core/n3515_172 ),
	.F(\top/processor/sha_core/n3515_148 )
);
defparam \top/processor/sha_core/n3515_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [4]),
	.I2(\top/processor/sha_core/w[1] [4]),
	.F(\top/processor/sha_core/n3515_149 )
);
defparam \top/processor/sha_core/n3515_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [4]),
	.I2(\top/processor/sha_core/w[5] [4]),
	.F(\top/processor/sha_core/n3515_150 )
);
defparam \top/processor/sha_core/n3515_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_172 ),
	.I3(\top/processor/sha_core/n3515_149 ),
	.F(\top/processor/sha_core/n3887_116 )
);
defparam \top/processor/sha_core/n3887_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [4]),
	.I2(\top/processor/sha_core/w[7] [4]),
	.F(\top/processor/sha_core/n3887_117 )
);
defparam \top/processor/sha_core/n3887_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_119 ),
	.I3(\top/processor/sha_core/n3515_173 ),
	.F(\top/processor/sha_core/n3515_151 )
);
defparam \top/processor/sha_core/n3515_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [4]),
	.I2(\top/processor/sha_core/w[9] [4]),
	.F(\top/processor/sha_core/n3515_152 )
);
defparam \top/processor/sha_core/n3515_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [4]),
	.I2(\top/processor/sha_core/w[13] [4]),
	.F(\top/processor/sha_core/n3515_153 )
);
defparam \top/processor/sha_core/n3515_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_173 ),
	.I3(\top/processor/sha_core/n3515_152 ),
	.F(\top/processor/sha_core/n3887_118 )
);
defparam \top/processor/sha_core/n3887_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [4]),
	.I2(\top/processor/sha_core/w[15] [4]),
	.F(\top/processor/sha_core/n3887_119 )
);
defparam \top/processor/sha_core/n3887_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_121 ),
	.I3(\top/processor/sha_core/n3515_174 ),
	.F(\top/processor/sha_core/n3515_154 )
);
defparam \top/processor/sha_core/n3515_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [4]),
	.I2(\top/processor/sha_core/w[17] [4]),
	.F(\top/processor/sha_core/n3515_155 )
);
defparam \top/processor/sha_core/n3515_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [4]),
	.I2(\top/processor/sha_core/w[21] [4]),
	.F(\top/processor/sha_core/n3515_156 )
);
defparam \top/processor/sha_core/n3515_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_174 ),
	.I3(\top/processor/sha_core/n3515_155 ),
	.F(\top/processor/sha_core/n3887_120 )
);
defparam \top/processor/sha_core/n3887_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [4]),
	.I2(\top/processor/sha_core/w[23] [4]),
	.F(\top/processor/sha_core/n3887_121 )
);
defparam \top/processor/sha_core/n3887_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_123 ),
	.I3(\top/processor/sha_core/n3515_175 ),
	.F(\top/processor/sha_core/n3515_157 )
);
defparam \top/processor/sha_core/n3515_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [4]),
	.I2(\top/processor/sha_core/w[25] [4]),
	.F(\top/processor/sha_core/n3515_158 )
);
defparam \top/processor/sha_core/n3515_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [4]),
	.I2(\top/processor/sha_core/w[29] [4]),
	.F(\top/processor/sha_core/n3515_159 )
);
defparam \top/processor/sha_core/n3515_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_175 ),
	.I3(\top/processor/sha_core/n3515_158 ),
	.F(\top/processor/sha_core/n3887_122 )
);
defparam \top/processor/sha_core/n3887_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [4]),
	.I2(\top/processor/sha_core/w[31] [4]),
	.F(\top/processor/sha_core/n3887_123 )
);
defparam \top/processor/sha_core/n3887_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_127 ),
	.I3(\top/processor/sha_core/n3490_177 ),
	.F(\top/processor/sha_core/n3490_163 )
);
defparam \top/processor/sha_core/n3490_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [29]),
	.I2(\top/processor/sha_core/w[41] [29]),
	.F(\top/processor/sha_core/n3490_164 )
);
defparam \top/processor/sha_core/n3490_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [29]),
	.I2(\top/processor/sha_core/w[45] [29]),
	.F(\top/processor/sha_core/n3490_165 )
);
defparam \top/processor/sha_core/n3490_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_177 ),
	.I3(\top/processor/sha_core/n3490_164 ),
	.F(\top/processor/sha_core/n3862_126 )
);
defparam \top/processor/sha_core/n3862_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [29]),
	.I2(\top/processor/sha_core/w[47] [29]),
	.F(\top/processor/sha_core/n3862_127 )
);
defparam \top/processor/sha_core/n3862_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_125 ),
	.I3(\top/processor/sha_core/n3515_176 ),
	.F(\top/processor/sha_core/n3515_160 )
);
defparam \top/processor/sha_core/n3515_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [4]),
	.I2(\top/processor/sha_core/w[33] [4]),
	.F(\top/processor/sha_core/n3515_161 )
);
defparam \top/processor/sha_core/n3515_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [4]),
	.I2(\top/processor/sha_core/w[37] [4]),
	.F(\top/processor/sha_core/n3515_162 )
);
defparam \top/processor/sha_core/n3515_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_176 ),
	.I3(\top/processor/sha_core/n3515_161 ),
	.F(\top/processor/sha_core/n3887_124 )
);
defparam \top/processor/sha_core/n3887_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [4]),
	.I2(\top/processor/sha_core/w[39] [4]),
	.F(\top/processor/sha_core/n3887_125 )
);
defparam \top/processor/sha_core/n3887_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_127 ),
	.I3(\top/processor/sha_core/n3515_177 ),
	.F(\top/processor/sha_core/n3515_163 )
);
defparam \top/processor/sha_core/n3515_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [4]),
	.I2(\top/processor/sha_core/w[41] [4]),
	.F(\top/processor/sha_core/n3515_164 )
);
defparam \top/processor/sha_core/n3515_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [4]),
	.I2(\top/processor/sha_core/w[45] [4]),
	.F(\top/processor/sha_core/n3515_165 )
);
defparam \top/processor/sha_core/n3515_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_177 ),
	.I3(\top/processor/sha_core/n3515_164 ),
	.F(\top/processor/sha_core/n3887_126 )
);
defparam \top/processor/sha_core/n3887_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [4]),
	.I2(\top/processor/sha_core/w[47] [4]),
	.F(\top/processor/sha_core/n3887_127 )
);
defparam \top/processor/sha_core/n3887_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_129 ),
	.I3(\top/processor/sha_core/n3515_178 ),
	.F(\top/processor/sha_core/n3515_166 )
);
defparam \top/processor/sha_core/n3515_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [4]),
	.I2(\top/processor/sha_core/w[49] [4]),
	.F(\top/processor/sha_core/n3515_167 )
);
defparam \top/processor/sha_core/n3515_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [4]),
	.I2(\top/processor/sha_core/w[53] [4]),
	.F(\top/processor/sha_core/n3515_168 )
);
defparam \top/processor/sha_core/n3515_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_178 ),
	.I3(\top/processor/sha_core/n3515_167 ),
	.F(\top/processor/sha_core/n3887_128 )
);
defparam \top/processor/sha_core/n3887_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [4]),
	.I2(\top/processor/sha_core/w[55] [4]),
	.F(\top/processor/sha_core/n3887_129 )
);
defparam \top/processor/sha_core/n3887_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3515_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3887_131 ),
	.I3(\top/processor/sha_core/n3515_179 ),
	.F(\top/processor/sha_core/n3515_169 )
);
defparam \top/processor/sha_core/n3515_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3515_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [4]),
	.I2(\top/processor/sha_core/w[57] [4]),
	.F(\top/processor/sha_core/n3515_170 )
);
defparam \top/processor/sha_core/n3515_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [4]),
	.I2(\top/processor/sha_core/w[61] [4]),
	.F(\top/processor/sha_core/n3515_171 )
);
defparam \top/processor/sha_core/n3515_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3887_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3515_179 ),
	.I3(\top/processor/sha_core/n3515_170 ),
	.F(\top/processor/sha_core/n3887_130 )
);
defparam \top/processor/sha_core/n3887_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3887_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [4]),
	.I2(\top/processor/sha_core/w[63] [4]),
	.F(\top/processor/sha_core/n3887_131 )
);
defparam \top/processor/sha_core/n3887_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_117 ),
	.I3(\top/processor/sha_core/n3516_172 ),
	.F(\top/processor/sha_core/n3516_148 )
);
defparam \top/processor/sha_core/n3516_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [3]),
	.I2(\top/processor/sha_core/w[1] [3]),
	.F(\top/processor/sha_core/n3516_149 )
);
defparam \top/processor/sha_core/n3516_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [3]),
	.I2(\top/processor/sha_core/w[5] [3]),
	.F(\top/processor/sha_core/n3516_150 )
);
defparam \top/processor/sha_core/n3516_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_172 ),
	.I3(\top/processor/sha_core/n3516_149 ),
	.F(\top/processor/sha_core/n3888_116 )
);
defparam \top/processor/sha_core/n3888_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [3]),
	.I2(\top/processor/sha_core/w[7] [3]),
	.F(\top/processor/sha_core/n3888_117 )
);
defparam \top/processor/sha_core/n3888_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_119 ),
	.I3(\top/processor/sha_core/n3516_173 ),
	.F(\top/processor/sha_core/n3516_151 )
);
defparam \top/processor/sha_core/n3516_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [3]),
	.I2(\top/processor/sha_core/w[9] [3]),
	.F(\top/processor/sha_core/n3516_152 )
);
defparam \top/processor/sha_core/n3516_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [3]),
	.I2(\top/processor/sha_core/w[13] [3]),
	.F(\top/processor/sha_core/n3516_153 )
);
defparam \top/processor/sha_core/n3516_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_173 ),
	.I3(\top/processor/sha_core/n3516_152 ),
	.F(\top/processor/sha_core/n3888_118 )
);
defparam \top/processor/sha_core/n3888_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [3]),
	.I2(\top/processor/sha_core/w[15] [3]),
	.F(\top/processor/sha_core/n3888_119 )
);
defparam \top/processor/sha_core/n3888_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_121 ),
	.I3(\top/processor/sha_core/n3516_174 ),
	.F(\top/processor/sha_core/n3516_154 )
);
defparam \top/processor/sha_core/n3516_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [3]),
	.I2(\top/processor/sha_core/w[17] [3]),
	.F(\top/processor/sha_core/n3516_155 )
);
defparam \top/processor/sha_core/n3516_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [3]),
	.I2(\top/processor/sha_core/w[21] [3]),
	.F(\top/processor/sha_core/n3516_156 )
);
defparam \top/processor/sha_core/n3516_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_174 ),
	.I3(\top/processor/sha_core/n3516_155 ),
	.F(\top/processor/sha_core/n3888_120 )
);
defparam \top/processor/sha_core/n3888_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [3]),
	.I2(\top/processor/sha_core/w[23] [3]),
	.F(\top/processor/sha_core/n3888_121 )
);
defparam \top/processor/sha_core/n3888_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_123 ),
	.I3(\top/processor/sha_core/n3516_175 ),
	.F(\top/processor/sha_core/n3516_157 )
);
defparam \top/processor/sha_core/n3516_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [3]),
	.I2(\top/processor/sha_core/w[25] [3]),
	.F(\top/processor/sha_core/n3516_158 )
);
defparam \top/processor/sha_core/n3516_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [3]),
	.I2(\top/processor/sha_core/w[29] [3]),
	.F(\top/processor/sha_core/n3516_159 )
);
defparam \top/processor/sha_core/n3516_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_175 ),
	.I3(\top/processor/sha_core/n3516_158 ),
	.F(\top/processor/sha_core/n3888_122 )
);
defparam \top/processor/sha_core/n3888_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [3]),
	.I2(\top/processor/sha_core/w[31] [3]),
	.F(\top/processor/sha_core/n3888_123 )
);
defparam \top/processor/sha_core/n3888_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_125 ),
	.I3(\top/processor/sha_core/n3516_176 ),
	.F(\top/processor/sha_core/n3516_160 )
);
defparam \top/processor/sha_core/n3516_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [3]),
	.I2(\top/processor/sha_core/w[33] [3]),
	.F(\top/processor/sha_core/n3516_161 )
);
defparam \top/processor/sha_core/n3516_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [3]),
	.I2(\top/processor/sha_core/w[37] [3]),
	.F(\top/processor/sha_core/n3516_162 )
);
defparam \top/processor/sha_core/n3516_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_176 ),
	.I3(\top/processor/sha_core/n3516_161 ),
	.F(\top/processor/sha_core/n3888_124 )
);
defparam \top/processor/sha_core/n3888_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [3]),
	.I2(\top/processor/sha_core/w[39] [3]),
	.F(\top/processor/sha_core/n3888_125 )
);
defparam \top/processor/sha_core/n3888_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_127 ),
	.I3(\top/processor/sha_core/n3516_177 ),
	.F(\top/processor/sha_core/n3516_163 )
);
defparam \top/processor/sha_core/n3516_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [3]),
	.I2(\top/processor/sha_core/w[41] [3]),
	.F(\top/processor/sha_core/n3516_164 )
);
defparam \top/processor/sha_core/n3516_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [3]),
	.I2(\top/processor/sha_core/w[45] [3]),
	.F(\top/processor/sha_core/n3516_165 )
);
defparam \top/processor/sha_core/n3516_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_177 ),
	.I3(\top/processor/sha_core/n3516_164 ),
	.F(\top/processor/sha_core/n3888_126 )
);
defparam \top/processor/sha_core/n3888_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [3]),
	.I2(\top/processor/sha_core/w[47] [3]),
	.F(\top/processor/sha_core/n3888_127 )
);
defparam \top/processor/sha_core/n3888_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_129 ),
	.I3(\top/processor/sha_core/n3490_178 ),
	.F(\top/processor/sha_core/n3490_166 )
);
defparam \top/processor/sha_core/n3490_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [29]),
	.I2(\top/processor/sha_core/w[49] [29]),
	.F(\top/processor/sha_core/n3490_167 )
);
defparam \top/processor/sha_core/n3490_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [29]),
	.I2(\top/processor/sha_core/w[53] [29]),
	.F(\top/processor/sha_core/n3490_168 )
);
defparam \top/processor/sha_core/n3490_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_178 ),
	.I3(\top/processor/sha_core/n3490_167 ),
	.F(\top/processor/sha_core/n3862_128 )
);
defparam \top/processor/sha_core/n3862_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [29]),
	.I2(\top/processor/sha_core/w[55] [29]),
	.F(\top/processor/sha_core/n3862_129 )
);
defparam \top/processor/sha_core/n3862_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_129 ),
	.I3(\top/processor/sha_core/n3516_178 ),
	.F(\top/processor/sha_core/n3516_166 )
);
defparam \top/processor/sha_core/n3516_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [3]),
	.I2(\top/processor/sha_core/w[49] [3]),
	.F(\top/processor/sha_core/n3516_167 )
);
defparam \top/processor/sha_core/n3516_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [3]),
	.I2(\top/processor/sha_core/w[53] [3]),
	.F(\top/processor/sha_core/n3516_168 )
);
defparam \top/processor/sha_core/n3516_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_178 ),
	.I3(\top/processor/sha_core/n3516_167 ),
	.F(\top/processor/sha_core/n3888_128 )
);
defparam \top/processor/sha_core/n3888_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [3]),
	.I2(\top/processor/sha_core/w[55] [3]),
	.F(\top/processor/sha_core/n3888_129 )
);
defparam \top/processor/sha_core/n3888_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3516_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3888_131 ),
	.I3(\top/processor/sha_core/n3516_179 ),
	.F(\top/processor/sha_core/n3516_169 )
);
defparam \top/processor/sha_core/n3516_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3516_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [3]),
	.I2(\top/processor/sha_core/w[57] [3]),
	.F(\top/processor/sha_core/n3516_170 )
);
defparam \top/processor/sha_core/n3516_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [3]),
	.I2(\top/processor/sha_core/w[61] [3]),
	.F(\top/processor/sha_core/n3516_171 )
);
defparam \top/processor/sha_core/n3516_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3888_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3516_179 ),
	.I3(\top/processor/sha_core/n3516_170 ),
	.F(\top/processor/sha_core/n3888_130 )
);
defparam \top/processor/sha_core/n3888_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3888_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [3]),
	.I2(\top/processor/sha_core/w[63] [3]),
	.F(\top/processor/sha_core/n3888_131 )
);
defparam \top/processor/sha_core/n3888_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_117 ),
	.I3(\top/processor/sha_core/n3517_172 ),
	.F(\top/processor/sha_core/n3517_148 )
);
defparam \top/processor/sha_core/n3517_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [2]),
	.I2(\top/processor/sha_core/w[1] [2]),
	.F(\top/processor/sha_core/n3517_149 )
);
defparam \top/processor/sha_core/n3517_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [2]),
	.I2(\top/processor/sha_core/w[5] [2]),
	.F(\top/processor/sha_core/n3517_150 )
);
defparam \top/processor/sha_core/n3517_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_172 ),
	.I3(\top/processor/sha_core/n3517_149 ),
	.F(\top/processor/sha_core/n3889_116 )
);
defparam \top/processor/sha_core/n3889_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [2]),
	.I2(\top/processor/sha_core/w[7] [2]),
	.F(\top/processor/sha_core/n3889_117 )
);
defparam \top/processor/sha_core/n3889_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_119 ),
	.I3(\top/processor/sha_core/n3517_173 ),
	.F(\top/processor/sha_core/n3517_151 )
);
defparam \top/processor/sha_core/n3517_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [2]),
	.I2(\top/processor/sha_core/w[9] [2]),
	.F(\top/processor/sha_core/n3517_152 )
);
defparam \top/processor/sha_core/n3517_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [2]),
	.I2(\top/processor/sha_core/w[13] [2]),
	.F(\top/processor/sha_core/n3517_153 )
);
defparam \top/processor/sha_core/n3517_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_173 ),
	.I3(\top/processor/sha_core/n3517_152 ),
	.F(\top/processor/sha_core/n3889_118 )
);
defparam \top/processor/sha_core/n3889_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [2]),
	.I2(\top/processor/sha_core/w[15] [2]),
	.F(\top/processor/sha_core/n3889_119 )
);
defparam \top/processor/sha_core/n3889_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_121 ),
	.I3(\top/processor/sha_core/n3517_174 ),
	.F(\top/processor/sha_core/n3517_154 )
);
defparam \top/processor/sha_core/n3517_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [2]),
	.I2(\top/processor/sha_core/w[17] [2]),
	.F(\top/processor/sha_core/n3517_155 )
);
defparam \top/processor/sha_core/n3517_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [2]),
	.I2(\top/processor/sha_core/w[21] [2]),
	.F(\top/processor/sha_core/n3517_156 )
);
defparam \top/processor/sha_core/n3517_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_174 ),
	.I3(\top/processor/sha_core/n3517_155 ),
	.F(\top/processor/sha_core/n3889_120 )
);
defparam \top/processor/sha_core/n3889_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [2]),
	.I2(\top/processor/sha_core/w[23] [2]),
	.F(\top/processor/sha_core/n3889_121 )
);
defparam \top/processor/sha_core/n3889_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_123 ),
	.I3(\top/processor/sha_core/n3517_175 ),
	.F(\top/processor/sha_core/n3517_157 )
);
defparam \top/processor/sha_core/n3517_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [2]),
	.I2(\top/processor/sha_core/w[25] [2]),
	.F(\top/processor/sha_core/n3517_158 )
);
defparam \top/processor/sha_core/n3517_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [2]),
	.I2(\top/processor/sha_core/w[29] [2]),
	.F(\top/processor/sha_core/n3517_159 )
);
defparam \top/processor/sha_core/n3517_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_175 ),
	.I3(\top/processor/sha_core/n3517_158 ),
	.F(\top/processor/sha_core/n3889_122 )
);
defparam \top/processor/sha_core/n3889_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [2]),
	.I2(\top/processor/sha_core/w[31] [2]),
	.F(\top/processor/sha_core/n3889_123 )
);
defparam \top/processor/sha_core/n3889_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_125 ),
	.I3(\top/processor/sha_core/n3517_176 ),
	.F(\top/processor/sha_core/n3517_160 )
);
defparam \top/processor/sha_core/n3517_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [2]),
	.I2(\top/processor/sha_core/w[33] [2]),
	.F(\top/processor/sha_core/n3517_161 )
);
defparam \top/processor/sha_core/n3517_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [2]),
	.I2(\top/processor/sha_core/w[37] [2]),
	.F(\top/processor/sha_core/n3517_162 )
);
defparam \top/processor/sha_core/n3517_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_176 ),
	.I3(\top/processor/sha_core/n3517_161 ),
	.F(\top/processor/sha_core/n3889_124 )
);
defparam \top/processor/sha_core/n3889_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [2]),
	.I2(\top/processor/sha_core/w[39] [2]),
	.F(\top/processor/sha_core/n3889_125 )
);
defparam \top/processor/sha_core/n3889_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_127 ),
	.I3(\top/processor/sha_core/n3517_177 ),
	.F(\top/processor/sha_core/n3517_163 )
);
defparam \top/processor/sha_core/n3517_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [2]),
	.I2(\top/processor/sha_core/w[41] [2]),
	.F(\top/processor/sha_core/n3517_164 )
);
defparam \top/processor/sha_core/n3517_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [2]),
	.I2(\top/processor/sha_core/w[45] [2]),
	.F(\top/processor/sha_core/n3517_165 )
);
defparam \top/processor/sha_core/n3517_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_177 ),
	.I3(\top/processor/sha_core/n3517_164 ),
	.F(\top/processor/sha_core/n3889_126 )
);
defparam \top/processor/sha_core/n3889_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [2]),
	.I2(\top/processor/sha_core/w[47] [2]),
	.F(\top/processor/sha_core/n3889_127 )
);
defparam \top/processor/sha_core/n3889_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_129 ),
	.I3(\top/processor/sha_core/n3517_178 ),
	.F(\top/processor/sha_core/n3517_166 )
);
defparam \top/processor/sha_core/n3517_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [2]),
	.I2(\top/processor/sha_core/w[49] [2]),
	.F(\top/processor/sha_core/n3517_167 )
);
defparam \top/processor/sha_core/n3517_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [2]),
	.I2(\top/processor/sha_core/w[53] [2]),
	.F(\top/processor/sha_core/n3517_168 )
);
defparam \top/processor/sha_core/n3517_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_178 ),
	.I3(\top/processor/sha_core/n3517_167 ),
	.F(\top/processor/sha_core/n3889_128 )
);
defparam \top/processor/sha_core/n3889_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [2]),
	.I2(\top/processor/sha_core/w[55] [2]),
	.F(\top/processor/sha_core/n3889_129 )
);
defparam \top/processor/sha_core/n3889_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3517_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3889_131 ),
	.I3(\top/processor/sha_core/n3517_179 ),
	.F(\top/processor/sha_core/n3517_169 )
);
defparam \top/processor/sha_core/n3517_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3517_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [2]),
	.I2(\top/processor/sha_core/w[57] [2]),
	.F(\top/processor/sha_core/n3517_170 )
);
defparam \top/processor/sha_core/n3517_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [2]),
	.I2(\top/processor/sha_core/w[61] [2]),
	.F(\top/processor/sha_core/n3517_171 )
);
defparam \top/processor/sha_core/n3517_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3889_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3517_179 ),
	.I3(\top/processor/sha_core/n3517_170 ),
	.F(\top/processor/sha_core/n3889_130 )
);
defparam \top/processor/sha_core/n3889_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3889_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [2]),
	.I2(\top/processor/sha_core/w[63] [2]),
	.F(\top/processor/sha_core/n3889_131 )
);
defparam \top/processor/sha_core/n3889_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3490_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3862_131 ),
	.I3(\top/processor/sha_core/n3490_179 ),
	.F(\top/processor/sha_core/n3490_169 )
);
defparam \top/processor/sha_core/n3490_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3490_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [29]),
	.I2(\top/processor/sha_core/w[57] [29]),
	.F(\top/processor/sha_core/n3490_170 )
);
defparam \top/processor/sha_core/n3490_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [29]),
	.I2(\top/processor/sha_core/w[61] [29]),
	.F(\top/processor/sha_core/n3490_171 )
);
defparam \top/processor/sha_core/n3490_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3862_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3490_179 ),
	.I3(\top/processor/sha_core/n3490_170 ),
	.F(\top/processor/sha_core/n3862_130 )
);
defparam \top/processor/sha_core/n3862_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3862_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [29]),
	.I2(\top/processor/sha_core/w[63] [29]),
	.F(\top/processor/sha_core/n3862_131 )
);
defparam \top/processor/sha_core/n3862_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_117 ),
	.I3(\top/processor/sha_core/n3518_172 ),
	.F(\top/processor/sha_core/n3518_148 )
);
defparam \top/processor/sha_core/n3518_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [1]),
	.I2(\top/processor/sha_core/w[1] [1]),
	.F(\top/processor/sha_core/n3518_149 )
);
defparam \top/processor/sha_core/n3518_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [1]),
	.I2(\top/processor/sha_core/w[5] [1]),
	.F(\top/processor/sha_core/n3518_150 )
);
defparam \top/processor/sha_core/n3518_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_172 ),
	.I3(\top/processor/sha_core/n3518_149 ),
	.F(\top/processor/sha_core/n3890_116 )
);
defparam \top/processor/sha_core/n3890_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [1]),
	.I2(\top/processor/sha_core/w[7] [1]),
	.F(\top/processor/sha_core/n3890_117 )
);
defparam \top/processor/sha_core/n3890_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_119 ),
	.I3(\top/processor/sha_core/n3518_173 ),
	.F(\top/processor/sha_core/n3518_151 )
);
defparam \top/processor/sha_core/n3518_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [1]),
	.I2(\top/processor/sha_core/w[9] [1]),
	.F(\top/processor/sha_core/n3518_152 )
);
defparam \top/processor/sha_core/n3518_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [1]),
	.I2(\top/processor/sha_core/w[13] [1]),
	.F(\top/processor/sha_core/n3518_153 )
);
defparam \top/processor/sha_core/n3518_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_173 ),
	.I3(\top/processor/sha_core/n3518_152 ),
	.F(\top/processor/sha_core/n3890_118 )
);
defparam \top/processor/sha_core/n3890_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [1]),
	.I2(\top/processor/sha_core/w[15] [1]),
	.F(\top/processor/sha_core/n3890_119 )
);
defparam \top/processor/sha_core/n3890_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_121 ),
	.I3(\top/processor/sha_core/n3518_174 ),
	.F(\top/processor/sha_core/n3518_154 )
);
defparam \top/processor/sha_core/n3518_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [1]),
	.I2(\top/processor/sha_core/w[17] [1]),
	.F(\top/processor/sha_core/n3518_155 )
);
defparam \top/processor/sha_core/n3518_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [1]),
	.I2(\top/processor/sha_core/w[21] [1]),
	.F(\top/processor/sha_core/n3518_156 )
);
defparam \top/processor/sha_core/n3518_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_174 ),
	.I3(\top/processor/sha_core/n3518_155 ),
	.F(\top/processor/sha_core/n3890_120 )
);
defparam \top/processor/sha_core/n3890_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [1]),
	.I2(\top/processor/sha_core/w[23] [1]),
	.F(\top/processor/sha_core/n3890_121 )
);
defparam \top/processor/sha_core/n3890_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_123 ),
	.I3(\top/processor/sha_core/n3518_175 ),
	.F(\top/processor/sha_core/n3518_157 )
);
defparam \top/processor/sha_core/n3518_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [1]),
	.I2(\top/processor/sha_core/w[25] [1]),
	.F(\top/processor/sha_core/n3518_158 )
);
defparam \top/processor/sha_core/n3518_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [1]),
	.I2(\top/processor/sha_core/w[29] [1]),
	.F(\top/processor/sha_core/n3518_159 )
);
defparam \top/processor/sha_core/n3518_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_175 ),
	.I3(\top/processor/sha_core/n3518_158 ),
	.F(\top/processor/sha_core/n3890_122 )
);
defparam \top/processor/sha_core/n3890_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [1]),
	.I2(\top/processor/sha_core/w[31] [1]),
	.F(\top/processor/sha_core/n3890_123 )
);
defparam \top/processor/sha_core/n3890_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_125 ),
	.I3(\top/processor/sha_core/n3518_176 ),
	.F(\top/processor/sha_core/n3518_160 )
);
defparam \top/processor/sha_core/n3518_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [1]),
	.I2(\top/processor/sha_core/w[33] [1]),
	.F(\top/processor/sha_core/n3518_161 )
);
defparam \top/processor/sha_core/n3518_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [1]),
	.I2(\top/processor/sha_core/w[37] [1]),
	.F(\top/processor/sha_core/n3518_162 )
);
defparam \top/processor/sha_core/n3518_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_176 ),
	.I3(\top/processor/sha_core/n3518_161 ),
	.F(\top/processor/sha_core/n3890_124 )
);
defparam \top/processor/sha_core/n3890_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [1]),
	.I2(\top/processor/sha_core/w[39] [1]),
	.F(\top/processor/sha_core/n3890_125 )
);
defparam \top/processor/sha_core/n3890_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_127 ),
	.I3(\top/processor/sha_core/n3518_177 ),
	.F(\top/processor/sha_core/n3518_163 )
);
defparam \top/processor/sha_core/n3518_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [1]),
	.I2(\top/processor/sha_core/w[41] [1]),
	.F(\top/processor/sha_core/n3518_164 )
);
defparam \top/processor/sha_core/n3518_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [1]),
	.I2(\top/processor/sha_core/w[45] [1]),
	.F(\top/processor/sha_core/n3518_165 )
);
defparam \top/processor/sha_core/n3518_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_177 ),
	.I3(\top/processor/sha_core/n3518_164 ),
	.F(\top/processor/sha_core/n3890_126 )
);
defparam \top/processor/sha_core/n3890_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [1]),
	.I2(\top/processor/sha_core/w[47] [1]),
	.F(\top/processor/sha_core/n3890_127 )
);
defparam \top/processor/sha_core/n3890_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_129 ),
	.I3(\top/processor/sha_core/n3518_178 ),
	.F(\top/processor/sha_core/n3518_166 )
);
defparam \top/processor/sha_core/n3518_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [1]),
	.I2(\top/processor/sha_core/w[49] [1]),
	.F(\top/processor/sha_core/n3518_167 )
);
defparam \top/processor/sha_core/n3518_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [1]),
	.I2(\top/processor/sha_core/w[53] [1]),
	.F(\top/processor/sha_core/n3518_168 )
);
defparam \top/processor/sha_core/n3518_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_178 ),
	.I3(\top/processor/sha_core/n3518_167 ),
	.F(\top/processor/sha_core/n3890_128 )
);
defparam \top/processor/sha_core/n3890_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [1]),
	.I2(\top/processor/sha_core/w[55] [1]),
	.F(\top/processor/sha_core/n3890_129 )
);
defparam \top/processor/sha_core/n3890_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3518_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3890_131 ),
	.I3(\top/processor/sha_core/n3518_179 ),
	.F(\top/processor/sha_core/n3518_169 )
);
defparam \top/processor/sha_core/n3518_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3518_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [1]),
	.I2(\top/processor/sha_core/w[57] [1]),
	.F(\top/processor/sha_core/n3518_170 )
);
defparam \top/processor/sha_core/n3518_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [1]),
	.I2(\top/processor/sha_core/w[61] [1]),
	.F(\top/processor/sha_core/n3518_171 )
);
defparam \top/processor/sha_core/n3518_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3890_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3518_179 ),
	.I3(\top/processor/sha_core/n3518_170 ),
	.F(\top/processor/sha_core/n3890_130 )
);
defparam \top/processor/sha_core/n3890_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3890_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [1]),
	.I2(\top/processor/sha_core/w[63] [1]),
	.F(\top/processor/sha_core/n3890_131 )
);
defparam \top/processor/sha_core/n3890_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_117 ),
	.I3(\top/processor/sha_core/n3519_172 ),
	.F(\top/processor/sha_core/n3519_148 )
);
defparam \top/processor/sha_core/n3519_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [0]),
	.I2(\top/processor/sha_core/w[1] [0]),
	.F(\top/processor/sha_core/n3519_149 )
);
defparam \top/processor/sha_core/n3519_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [0]),
	.I2(\top/processor/sha_core/w[5] [0]),
	.F(\top/processor/sha_core/n3519_150 )
);
defparam \top/processor/sha_core/n3519_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_172 ),
	.I3(\top/processor/sha_core/n3519_149 ),
	.F(\top/processor/sha_core/n3891_116 )
);
defparam \top/processor/sha_core/n3891_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [0]),
	.I2(\top/processor/sha_core/w[7] [0]),
	.F(\top/processor/sha_core/n3891_117 )
);
defparam \top/processor/sha_core/n3891_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_119 ),
	.I3(\top/processor/sha_core/n3519_173 ),
	.F(\top/processor/sha_core/n3519_151 )
);
defparam \top/processor/sha_core/n3519_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [0]),
	.I2(\top/processor/sha_core/w[9] [0]),
	.F(\top/processor/sha_core/n3519_152 )
);
defparam \top/processor/sha_core/n3519_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [0]),
	.I2(\top/processor/sha_core/w[13] [0]),
	.F(\top/processor/sha_core/n3519_153 )
);
defparam \top/processor/sha_core/n3519_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_173 ),
	.I3(\top/processor/sha_core/n3519_152 ),
	.F(\top/processor/sha_core/n3891_118 )
);
defparam \top/processor/sha_core/n3891_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [0]),
	.I2(\top/processor/sha_core/w[15] [0]),
	.F(\top/processor/sha_core/n3891_119 )
);
defparam \top/processor/sha_core/n3891_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3491_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_117 ),
	.I3(\top/processor/sha_core/n3491_172 ),
	.F(\top/processor/sha_core/n3491_148 )
);
defparam \top/processor/sha_core/n3491_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [28]),
	.I2(\top/processor/sha_core/w[1] [28]),
	.F(\top/processor/sha_core/n3491_149 )
);
defparam \top/processor/sha_core/n3491_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [28]),
	.I2(\top/processor/sha_core/w[5] [28]),
	.F(\top/processor/sha_core/n3491_150 )
);
defparam \top/processor/sha_core/n3491_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_172 ),
	.I3(\top/processor/sha_core/n3491_149 ),
	.F(\top/processor/sha_core/n3863_116 )
);
defparam \top/processor/sha_core/n3863_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [28]),
	.I2(\top/processor/sha_core/w[7] [28]),
	.F(\top/processor/sha_core/n3863_117 )
);
defparam \top/processor/sha_core/n3863_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_121 ),
	.I3(\top/processor/sha_core/n3519_174 ),
	.F(\top/processor/sha_core/n3519_154 )
);
defparam \top/processor/sha_core/n3519_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [0]),
	.I2(\top/processor/sha_core/w[17] [0]),
	.F(\top/processor/sha_core/n3519_155 )
);
defparam \top/processor/sha_core/n3519_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [0]),
	.I2(\top/processor/sha_core/w[21] [0]),
	.F(\top/processor/sha_core/n3519_156 )
);
defparam \top/processor/sha_core/n3519_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_174 ),
	.I3(\top/processor/sha_core/n3519_155 ),
	.F(\top/processor/sha_core/n3891_120 )
);
defparam \top/processor/sha_core/n3891_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [0]),
	.I2(\top/processor/sha_core/w[23] [0]),
	.F(\top/processor/sha_core/n3891_121 )
);
defparam \top/processor/sha_core/n3891_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_123 ),
	.I3(\top/processor/sha_core/n3519_175 ),
	.F(\top/processor/sha_core/n3519_157 )
);
defparam \top/processor/sha_core/n3519_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [0]),
	.I2(\top/processor/sha_core/w[25] [0]),
	.F(\top/processor/sha_core/n3519_158 )
);
defparam \top/processor/sha_core/n3519_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [0]),
	.I2(\top/processor/sha_core/w[29] [0]),
	.F(\top/processor/sha_core/n3519_159 )
);
defparam \top/processor/sha_core/n3519_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_175 ),
	.I3(\top/processor/sha_core/n3519_158 ),
	.F(\top/processor/sha_core/n3891_122 )
);
defparam \top/processor/sha_core/n3891_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [0]),
	.I2(\top/processor/sha_core/w[31] [0]),
	.F(\top/processor/sha_core/n3891_123 )
);
defparam \top/processor/sha_core/n3891_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_125 ),
	.I3(\top/processor/sha_core/n3519_176 ),
	.F(\top/processor/sha_core/n3519_160 )
);
defparam \top/processor/sha_core/n3519_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [0]),
	.I2(\top/processor/sha_core/w[33] [0]),
	.F(\top/processor/sha_core/n3519_161 )
);
defparam \top/processor/sha_core/n3519_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [0]),
	.I2(\top/processor/sha_core/w[37] [0]),
	.F(\top/processor/sha_core/n3519_162 )
);
defparam \top/processor/sha_core/n3519_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_176 ),
	.I3(\top/processor/sha_core/n3519_161 ),
	.F(\top/processor/sha_core/n3891_124 )
);
defparam \top/processor/sha_core/n3891_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [0]),
	.I2(\top/processor/sha_core/w[39] [0]),
	.F(\top/processor/sha_core/n3891_125 )
);
defparam \top/processor/sha_core/n3891_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_127 ),
	.I3(\top/processor/sha_core/n3519_177 ),
	.F(\top/processor/sha_core/n3519_163 )
);
defparam \top/processor/sha_core/n3519_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [0]),
	.I2(\top/processor/sha_core/w[41] [0]),
	.F(\top/processor/sha_core/n3519_164 )
);
defparam \top/processor/sha_core/n3519_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [0]),
	.I2(\top/processor/sha_core/w[45] [0]),
	.F(\top/processor/sha_core/n3519_165 )
);
defparam \top/processor/sha_core/n3519_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_177 ),
	.I3(\top/processor/sha_core/n3519_164 ),
	.F(\top/processor/sha_core/n3891_126 )
);
defparam \top/processor/sha_core/n3891_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [0]),
	.I2(\top/processor/sha_core/w[47] [0]),
	.F(\top/processor/sha_core/n3891_127 )
);
defparam \top/processor/sha_core/n3891_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_129 ),
	.I3(\top/processor/sha_core/n3519_178 ),
	.F(\top/processor/sha_core/n3519_166 )
);
defparam \top/processor/sha_core/n3519_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [0]),
	.I2(\top/processor/sha_core/w[49] [0]),
	.F(\top/processor/sha_core/n3519_167 )
);
defparam \top/processor/sha_core/n3519_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [0]),
	.I2(\top/processor/sha_core/w[53] [0]),
	.F(\top/processor/sha_core/n3519_168 )
);
defparam \top/processor/sha_core/n3519_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_178 ),
	.I3(\top/processor/sha_core/n3519_167 ),
	.F(\top/processor/sha_core/n3891_128 )
);
defparam \top/processor/sha_core/n3891_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [0]),
	.I2(\top/processor/sha_core/w[55] [0]),
	.F(\top/processor/sha_core/n3891_129 )
);
defparam \top/processor/sha_core/n3891_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3519_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3891_131 ),
	.I3(\top/processor/sha_core/n3519_179 ),
	.F(\top/processor/sha_core/n3519_169 )
);
defparam \top/processor/sha_core/n3519_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3519_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [0]),
	.I2(\top/processor/sha_core/w[57] [0]),
	.F(\top/processor/sha_core/n3519_170 )
);
defparam \top/processor/sha_core/n3519_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [0]),
	.I2(\top/processor/sha_core/w[61] [0]),
	.F(\top/processor/sha_core/n3519_171 )
);
defparam \top/processor/sha_core/n3519_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3891_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3519_179 ),
	.I3(\top/processor/sha_core/n3519_170 ),
	.F(\top/processor/sha_core/n3891_130 )
);
defparam \top/processor/sha_core/n3891_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3891_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [0]),
	.I2(\top/processor/sha_core/w[63] [0]),
	.F(\top/processor/sha_core/n3891_131 )
);
defparam \top/processor/sha_core/n3891_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [31]),
	.I3(\top/processor/sha_core/w[1] [31]),
	.F(\top/processor/sha_core/n3607_172 )
);
defparam \top/processor/sha_core/n3607_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [30]),
	.I3(\top/processor/sha_core/w[1] [30]),
	.F(\top/processor/sha_core/n3608_172 )
);
defparam \top/processor/sha_core/n3608_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [29]),
	.I3(\top/processor/sha_core/w[1] [29]),
	.F(\top/processor/sha_core/n3609_172 )
);
defparam \top/processor/sha_core/n3609_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [28]),
	.I3(\top/processor/sha_core/w[1] [28]),
	.F(\top/processor/sha_core/n3610_172 )
);
defparam \top/processor/sha_core/n3610_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [27]),
	.I3(\top/processor/sha_core/w[1] [27]),
	.F(\top/processor/sha_core/n3611_172 )
);
defparam \top/processor/sha_core/n3611_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [26]),
	.I3(\top/processor/sha_core/w[1] [26]),
	.F(\top/processor/sha_core/n3612_172 )
);
defparam \top/processor/sha_core/n3612_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [25]),
	.I3(\top/processor/sha_core/w[1] [25]),
	.F(\top/processor/sha_core/n3613_172 )
);
defparam \top/processor/sha_core/n3613_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3491_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_119 ),
	.I3(\top/processor/sha_core/n3491_173 ),
	.F(\top/processor/sha_core/n3491_151 )
);
defparam \top/processor/sha_core/n3491_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [28]),
	.I2(\top/processor/sha_core/w[9] [28]),
	.F(\top/processor/sha_core/n3491_152 )
);
defparam \top/processor/sha_core/n3491_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [28]),
	.I2(\top/processor/sha_core/w[13] [28]),
	.F(\top/processor/sha_core/n3491_153 )
);
defparam \top/processor/sha_core/n3491_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_173 ),
	.I3(\top/processor/sha_core/n3491_152 ),
	.F(\top/processor/sha_core/n3863_118 )
);
defparam \top/processor/sha_core/n3863_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [28]),
	.I2(\top/processor/sha_core/w[15] [28]),
	.F(\top/processor/sha_core/n3863_119 )
);
defparam \top/processor/sha_core/n3863_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3614_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [24]),
	.I3(\top/processor/sha_core/w[1] [24]),
	.F(\top/processor/sha_core/n3614_172 )
);
defparam \top/processor/sha_core/n3614_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [23]),
	.I3(\top/processor/sha_core/w[1] [23]),
	.F(\top/processor/sha_core/n3615_172 )
);
defparam \top/processor/sha_core/n3615_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [22]),
	.I3(\top/processor/sha_core/w[1] [22]),
	.F(\top/processor/sha_core/n3616_172 )
);
defparam \top/processor/sha_core/n3616_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [21]),
	.I3(\top/processor/sha_core/w[1] [21]),
	.F(\top/processor/sha_core/n3617_172 )
);
defparam \top/processor/sha_core/n3617_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [20]),
	.I3(\top/processor/sha_core/w[1] [20]),
	.F(\top/processor/sha_core/n3618_172 )
);
defparam \top/processor/sha_core/n3618_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [19]),
	.I3(\top/processor/sha_core/w[1] [19]),
	.F(\top/processor/sha_core/n3619_172 )
);
defparam \top/processor/sha_core/n3619_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [18]),
	.I3(\top/processor/sha_core/w[1] [18]),
	.F(\top/processor/sha_core/n3620_172 )
);
defparam \top/processor/sha_core/n3620_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [17]),
	.I3(\top/processor/sha_core/w[1] [17]),
	.F(\top/processor/sha_core/n3621_172 )
);
defparam \top/processor/sha_core/n3621_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [16]),
	.I3(\top/processor/sha_core/w[1] [16]),
	.F(\top/processor/sha_core/n3622_172 )
);
defparam \top/processor/sha_core/n3622_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [15]),
	.I3(\top/processor/sha_core/w[1] [15]),
	.F(\top/processor/sha_core/n3623_172 )
);
defparam \top/processor/sha_core/n3623_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [14]),
	.I3(\top/processor/sha_core/w[1] [14]),
	.F(\top/processor/sha_core/n3624_172 )
);
defparam \top/processor/sha_core/n3624_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [13]),
	.I3(\top/processor/sha_core/w[1] [13]),
	.F(\top/processor/sha_core/n3625_172 )
);
defparam \top/processor/sha_core/n3625_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [12]),
	.I3(\top/processor/sha_core/w[1] [12]),
	.F(\top/processor/sha_core/n3626_172 )
);
defparam \top/processor/sha_core/n3626_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [11]),
	.I3(\top/processor/sha_core/w[1] [11]),
	.F(\top/processor/sha_core/n3627_172 )
);
defparam \top/processor/sha_core/n3627_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [10]),
	.I3(\top/processor/sha_core/w[1] [10]),
	.F(\top/processor/sha_core/n3628_172 )
);
defparam \top/processor/sha_core/n3628_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [9]),
	.I3(\top/processor/sha_core/w[1] [9]),
	.F(\top/processor/sha_core/n3629_172 )
);
defparam \top/processor/sha_core/n3629_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [8]),
	.I3(\top/processor/sha_core/w[1] [8]),
	.F(\top/processor/sha_core/n3630_172 )
);
defparam \top/processor/sha_core/n3630_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [7]),
	.I3(\top/processor/sha_core/w[1] [7]),
	.F(\top/processor/sha_core/n3631_172 )
);
defparam \top/processor/sha_core/n3631_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [6]),
	.I3(\top/processor/sha_core/w[1] [6]),
	.F(\top/processor/sha_core/n3632_172 )
);
defparam \top/processor/sha_core/n3632_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [5]),
	.I3(\top/processor/sha_core/w[1] [5]),
	.F(\top/processor/sha_core/n3633_172 )
);
defparam \top/processor/sha_core/n3633_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3491_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_121 ),
	.I3(\top/processor/sha_core/n3491_174 ),
	.F(\top/processor/sha_core/n3491_154 )
);
defparam \top/processor/sha_core/n3491_s141 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3491_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [28]),
	.I2(\top/processor/sha_core/w[17] [28]),
	.F(\top/processor/sha_core/n3491_155 )
);
defparam \top/processor/sha_core/n3491_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [28]),
	.I2(\top/processor/sha_core/w[21] [28]),
	.F(\top/processor/sha_core/n3491_156 )
);
defparam \top/processor/sha_core/n3491_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_174 ),
	.I3(\top/processor/sha_core/n3491_155 ),
	.F(\top/processor/sha_core/n3863_120 )
);
defparam \top/processor/sha_core/n3863_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [28]),
	.I2(\top/processor/sha_core/w[23] [28]),
	.F(\top/processor/sha_core/n3863_121 )
);
defparam \top/processor/sha_core/n3863_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3634_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [4]),
	.I3(\top/processor/sha_core/w[1] [4]),
	.F(\top/processor/sha_core/n3634_172 )
);
defparam \top/processor/sha_core/n3634_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [3]),
	.I3(\top/processor/sha_core/w[1] [3]),
	.F(\top/processor/sha_core/n3635_172 )
);
defparam \top/processor/sha_core/n3635_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [2]),
	.I3(\top/processor/sha_core/w[1] [2]),
	.F(\top/processor/sha_core/n3636_172 )
);
defparam \top/processor/sha_core/n3636_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [1]),
	.I3(\top/processor/sha_core/w[1] [1]),
	.F(\top/processor/sha_core/n3637_172 )
);
defparam \top/processor/sha_core/n3637_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[3] [0]),
	.I3(\top/processor/sha_core/w[1] [0]),
	.F(\top/processor/sha_core/n3638_172 )
);
defparam \top/processor/sha_core/n3638_s151 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3491_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_123 ),
	.I3(\top/processor/sha_core/n3491_175 ),
	.F(\top/processor/sha_core/n3491_157 )
);
defparam \top/processor/sha_core/n3491_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [28]),
	.I2(\top/processor/sha_core/w[25] [28]),
	.F(\top/processor/sha_core/n3491_158 )
);
defparam \top/processor/sha_core/n3491_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [28]),
	.I2(\top/processor/sha_core/w[29] [28]),
	.F(\top/processor/sha_core/n3491_159 )
);
defparam \top/processor/sha_core/n3491_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_175 ),
	.I3(\top/processor/sha_core/n3491_158 ),
	.F(\top/processor/sha_core/n3863_122 )
);
defparam \top/processor/sha_core/n3863_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [28]),
	.I2(\top/processor/sha_core/w[31] [28]),
	.F(\top/processor/sha_core/n3863_123 )
);
defparam \top/processor/sha_core/n3863_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [31]),
	.I3(\top/processor/sha_core/w[5] [31]),
	.F(\top/processor/sha_core/n3607_173 )
);
defparam \top/processor/sha_core/n3607_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [30]),
	.I3(\top/processor/sha_core/w[5] [30]),
	.F(\top/processor/sha_core/n3608_173 )
);
defparam \top/processor/sha_core/n3608_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [29]),
	.I3(\top/processor/sha_core/w[5] [29]),
	.F(\top/processor/sha_core/n3609_173 )
);
defparam \top/processor/sha_core/n3609_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3491_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_125 ),
	.I3(\top/processor/sha_core/n3491_176 ),
	.F(\top/processor/sha_core/n3491_160 )
);
defparam \top/processor/sha_core/n3491_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [28]),
	.I2(\top/processor/sha_core/w[33] [28]),
	.F(\top/processor/sha_core/n3491_161 )
);
defparam \top/processor/sha_core/n3491_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [28]),
	.I2(\top/processor/sha_core/w[37] [28]),
	.F(\top/processor/sha_core/n3491_162 )
);
defparam \top/processor/sha_core/n3491_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_176 ),
	.I3(\top/processor/sha_core/n3491_161 ),
	.F(\top/processor/sha_core/n3863_124 )
);
defparam \top/processor/sha_core/n3863_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [28]),
	.I2(\top/processor/sha_core/w[39] [28]),
	.F(\top/processor/sha_core/n3863_125 )
);
defparam \top/processor/sha_core/n3863_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3610_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [28]),
	.I3(\top/processor/sha_core/w[5] [28]),
	.F(\top/processor/sha_core/n3610_173 )
);
defparam \top/processor/sha_core/n3610_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [27]),
	.I3(\top/processor/sha_core/w[5] [27]),
	.F(\top/processor/sha_core/n3611_173 )
);
defparam \top/processor/sha_core/n3611_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [26]),
	.I3(\top/processor/sha_core/w[5] [26]),
	.F(\top/processor/sha_core/n3612_173 )
);
defparam \top/processor/sha_core/n3612_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [25]),
	.I3(\top/processor/sha_core/w[5] [25]),
	.F(\top/processor/sha_core/n3613_173 )
);
defparam \top/processor/sha_core/n3613_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [24]),
	.I3(\top/processor/sha_core/w[5] [24]),
	.F(\top/processor/sha_core/n3614_173 )
);
defparam \top/processor/sha_core/n3614_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [23]),
	.I3(\top/processor/sha_core/w[5] [23]),
	.F(\top/processor/sha_core/n3615_173 )
);
defparam \top/processor/sha_core/n3615_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [22]),
	.I3(\top/processor/sha_core/w[5] [22]),
	.F(\top/processor/sha_core/n3616_173 )
);
defparam \top/processor/sha_core/n3616_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [21]),
	.I3(\top/processor/sha_core/w[5] [21]),
	.F(\top/processor/sha_core/n3617_173 )
);
defparam \top/processor/sha_core/n3617_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [20]),
	.I3(\top/processor/sha_core/w[5] [20]),
	.F(\top/processor/sha_core/n3618_173 )
);
defparam \top/processor/sha_core/n3618_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [19]),
	.I3(\top/processor/sha_core/w[5] [19]),
	.F(\top/processor/sha_core/n3619_173 )
);
defparam \top/processor/sha_core/n3619_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [18]),
	.I3(\top/processor/sha_core/w[5] [18]),
	.F(\top/processor/sha_core/n3620_173 )
);
defparam \top/processor/sha_core/n3620_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [17]),
	.I3(\top/processor/sha_core/w[5] [17]),
	.F(\top/processor/sha_core/n3621_173 )
);
defparam \top/processor/sha_core/n3621_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [16]),
	.I3(\top/processor/sha_core/w[5] [16]),
	.F(\top/processor/sha_core/n3622_173 )
);
defparam \top/processor/sha_core/n3622_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [15]),
	.I3(\top/processor/sha_core/w[5] [15]),
	.F(\top/processor/sha_core/n3623_173 )
);
defparam \top/processor/sha_core/n3623_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [14]),
	.I3(\top/processor/sha_core/w[5] [14]),
	.F(\top/processor/sha_core/n3624_173 )
);
defparam \top/processor/sha_core/n3624_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [13]),
	.I3(\top/processor/sha_core/w[5] [13]),
	.F(\top/processor/sha_core/n3625_173 )
);
defparam \top/processor/sha_core/n3625_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [12]),
	.I3(\top/processor/sha_core/w[5] [12]),
	.F(\top/processor/sha_core/n3626_173 )
);
defparam \top/processor/sha_core/n3626_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [11]),
	.I3(\top/processor/sha_core/w[5] [11]),
	.F(\top/processor/sha_core/n3627_173 )
);
defparam \top/processor/sha_core/n3627_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [10]),
	.I3(\top/processor/sha_core/w[5] [10]),
	.F(\top/processor/sha_core/n3628_173 )
);
defparam \top/processor/sha_core/n3628_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [9]),
	.I3(\top/processor/sha_core/w[5] [9]),
	.F(\top/processor/sha_core/n3629_173 )
);
defparam \top/processor/sha_core/n3629_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3491_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_127 ),
	.I3(\top/processor/sha_core/n3491_177 ),
	.F(\top/processor/sha_core/n3491_163 )
);
defparam \top/processor/sha_core/n3491_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [28]),
	.I2(\top/processor/sha_core/w[41] [28]),
	.F(\top/processor/sha_core/n3491_164 )
);
defparam \top/processor/sha_core/n3491_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [28]),
	.I2(\top/processor/sha_core/w[45] [28]),
	.F(\top/processor/sha_core/n3491_165 )
);
defparam \top/processor/sha_core/n3491_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_177 ),
	.I3(\top/processor/sha_core/n3491_164 ),
	.F(\top/processor/sha_core/n3863_126 )
);
defparam \top/processor/sha_core/n3863_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [28]),
	.I2(\top/processor/sha_core/w[47] [28]),
	.F(\top/processor/sha_core/n3863_127 )
);
defparam \top/processor/sha_core/n3863_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_127 ),
	.I3(\top/processor/sha_core/n3488_177 ),
	.F(\top/processor/sha_core/n3488_163 )
);
defparam \top/processor/sha_core/n3488_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [31]),
	.I2(\top/processor/sha_core/w[17] [31]),
	.F(\top/processor/sha_core/n3488_164 )
);
defparam \top/processor/sha_core/n3488_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [31]),
	.I2(\top/processor/sha_core/w[21] [31]),
	.F(\top/processor/sha_core/n3488_165 )
);
defparam \top/processor/sha_core/n3488_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_177 ),
	.I3(\top/processor/sha_core/n3488_164 ),
	.F(\top/processor/sha_core/n3860_126 )
);
defparam \top/processor/sha_core/n3860_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [31]),
	.I2(\top/processor/sha_core/w[23] [31]),
	.F(\top/processor/sha_core/n3860_127 )
);
defparam \top/processor/sha_core/n3860_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3630_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [8]),
	.I3(\top/processor/sha_core/w[5] [8]),
	.F(\top/processor/sha_core/n3630_173 )
);
defparam \top/processor/sha_core/n3630_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [7]),
	.I3(\top/processor/sha_core/w[5] [7]),
	.F(\top/processor/sha_core/n3631_173 )
);
defparam \top/processor/sha_core/n3631_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [6]),
	.I3(\top/processor/sha_core/w[5] [6]),
	.F(\top/processor/sha_core/n3632_173 )
);
defparam \top/processor/sha_core/n3632_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [5]),
	.I3(\top/processor/sha_core/w[5] [5]),
	.F(\top/processor/sha_core/n3633_173 )
);
defparam \top/processor/sha_core/n3633_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [4]),
	.I3(\top/processor/sha_core/w[5] [4]),
	.F(\top/processor/sha_core/n3634_173 )
);
defparam \top/processor/sha_core/n3634_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [3]),
	.I3(\top/processor/sha_core/w[5] [3]),
	.F(\top/processor/sha_core/n3635_173 )
);
defparam \top/processor/sha_core/n3635_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [2]),
	.I3(\top/processor/sha_core/w[5] [2]),
	.F(\top/processor/sha_core/n3636_173 )
);
defparam \top/processor/sha_core/n3636_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [1]),
	.I3(\top/processor/sha_core/w[5] [1]),
	.F(\top/processor/sha_core/n3637_173 )
);
defparam \top/processor/sha_core/n3637_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[7] [0]),
	.I3(\top/processor/sha_core/w[5] [0]),
	.F(\top/processor/sha_core/n3638_173 )
);
defparam \top/processor/sha_core/n3638_s152 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3491_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_129 ),
	.I3(\top/processor/sha_core/n3491_178 ),
	.F(\top/processor/sha_core/n3491_166 )
);
defparam \top/processor/sha_core/n3491_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [28]),
	.I2(\top/processor/sha_core/w[49] [28]),
	.F(\top/processor/sha_core/n3491_167 )
);
defparam \top/processor/sha_core/n3491_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [28]),
	.I2(\top/processor/sha_core/w[53] [28]),
	.F(\top/processor/sha_core/n3491_168 )
);
defparam \top/processor/sha_core/n3491_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_178 ),
	.I3(\top/processor/sha_core/n3491_167 ),
	.F(\top/processor/sha_core/n3863_128 )
);
defparam \top/processor/sha_core/n3863_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [28]),
	.I2(\top/processor/sha_core/w[55] [28]),
	.F(\top/processor/sha_core/n3863_129 )
);
defparam \top/processor/sha_core/n3863_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3491_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3863_131 ),
	.I3(\top/processor/sha_core/n3491_179 ),
	.F(\top/processor/sha_core/n3491_169 )
);
defparam \top/processor/sha_core/n3491_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3491_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [28]),
	.I2(\top/processor/sha_core/w[57] [28]),
	.F(\top/processor/sha_core/n3491_170 )
);
defparam \top/processor/sha_core/n3491_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [28]),
	.I2(\top/processor/sha_core/w[61] [28]),
	.F(\top/processor/sha_core/n3491_171 )
);
defparam \top/processor/sha_core/n3491_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3863_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3491_179 ),
	.I3(\top/processor/sha_core/n3491_170 ),
	.F(\top/processor/sha_core/n3863_130 )
);
defparam \top/processor/sha_core/n3863_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3863_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [28]),
	.I2(\top/processor/sha_core/w[63] [28]),
	.F(\top/processor/sha_core/n3863_131 )
);
defparam \top/processor/sha_core/n3863_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [31]),
	.I3(\top/processor/sha_core/w[9] [31]),
	.F(\top/processor/sha_core/n3607_174 )
);
defparam \top/processor/sha_core/n3607_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [30]),
	.I3(\top/processor/sha_core/w[9] [30]),
	.F(\top/processor/sha_core/n3608_174 )
);
defparam \top/processor/sha_core/n3608_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [29]),
	.I3(\top/processor/sha_core/w[9] [29]),
	.F(\top/processor/sha_core/n3609_174 )
);
defparam \top/processor/sha_core/n3609_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [28]),
	.I3(\top/processor/sha_core/w[9] [28]),
	.F(\top/processor/sha_core/n3610_174 )
);
defparam \top/processor/sha_core/n3610_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [27]),
	.I3(\top/processor/sha_core/w[9] [27]),
	.F(\top/processor/sha_core/n3611_174 )
);
defparam \top/processor/sha_core/n3611_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [26]),
	.I3(\top/processor/sha_core/w[9] [26]),
	.F(\top/processor/sha_core/n3612_174 )
);
defparam \top/processor/sha_core/n3612_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [25]),
	.I3(\top/processor/sha_core/w[9] [25]),
	.F(\top/processor/sha_core/n3613_174 )
);
defparam \top/processor/sha_core/n3613_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [24]),
	.I3(\top/processor/sha_core/w[9] [24]),
	.F(\top/processor/sha_core/n3614_174 )
);
defparam \top/processor/sha_core/n3614_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [23]),
	.I3(\top/processor/sha_core/w[9] [23]),
	.F(\top/processor/sha_core/n3615_174 )
);
defparam \top/processor/sha_core/n3615_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [22]),
	.I3(\top/processor/sha_core/w[9] [22]),
	.F(\top/processor/sha_core/n3616_174 )
);
defparam \top/processor/sha_core/n3616_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [21]),
	.I3(\top/processor/sha_core/w[9] [21]),
	.F(\top/processor/sha_core/n3617_174 )
);
defparam \top/processor/sha_core/n3617_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [20]),
	.I3(\top/processor/sha_core/w[9] [20]),
	.F(\top/processor/sha_core/n3618_174 )
);
defparam \top/processor/sha_core/n3618_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [19]),
	.I3(\top/processor/sha_core/w[9] [19]),
	.F(\top/processor/sha_core/n3619_174 )
);
defparam \top/processor/sha_core/n3619_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [18]),
	.I3(\top/processor/sha_core/w[9] [18]),
	.F(\top/processor/sha_core/n3620_174 )
);
defparam \top/processor/sha_core/n3620_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [17]),
	.I3(\top/processor/sha_core/w[9] [17]),
	.F(\top/processor/sha_core/n3621_174 )
);
defparam \top/processor/sha_core/n3621_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [16]),
	.I3(\top/processor/sha_core/w[9] [16]),
	.F(\top/processor/sha_core/n3622_174 )
);
defparam \top/processor/sha_core/n3622_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [15]),
	.I3(\top/processor/sha_core/w[9] [15]),
	.F(\top/processor/sha_core/n3623_174 )
);
defparam \top/processor/sha_core/n3623_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [14]),
	.I3(\top/processor/sha_core/w[9] [14]),
	.F(\top/processor/sha_core/n3624_174 )
);
defparam \top/processor/sha_core/n3624_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [13]),
	.I3(\top/processor/sha_core/w[9] [13]),
	.F(\top/processor/sha_core/n3625_174 )
);
defparam \top/processor/sha_core/n3625_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3492_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_117 ),
	.I3(\top/processor/sha_core/n3492_172 ),
	.F(\top/processor/sha_core/n3492_148 )
);
defparam \top/processor/sha_core/n3492_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [27]),
	.I2(\top/processor/sha_core/w[1] [27]),
	.F(\top/processor/sha_core/n3492_149 )
);
defparam \top/processor/sha_core/n3492_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [27]),
	.I2(\top/processor/sha_core/w[5] [27]),
	.F(\top/processor/sha_core/n3492_150 )
);
defparam \top/processor/sha_core/n3492_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_172 ),
	.I3(\top/processor/sha_core/n3492_149 ),
	.F(\top/processor/sha_core/n3864_116 )
);
defparam \top/processor/sha_core/n3864_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [27]),
	.I2(\top/processor/sha_core/w[7] [27]),
	.F(\top/processor/sha_core/n3864_117 )
);
defparam \top/processor/sha_core/n3864_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3626_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [12]),
	.I3(\top/processor/sha_core/w[9] [12]),
	.F(\top/processor/sha_core/n3626_174 )
);
defparam \top/processor/sha_core/n3626_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [11]),
	.I3(\top/processor/sha_core/w[9] [11]),
	.F(\top/processor/sha_core/n3627_174 )
);
defparam \top/processor/sha_core/n3627_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [10]),
	.I3(\top/processor/sha_core/w[9] [10]),
	.F(\top/processor/sha_core/n3628_174 )
);
defparam \top/processor/sha_core/n3628_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [9]),
	.I3(\top/processor/sha_core/w[9] [9]),
	.F(\top/processor/sha_core/n3629_174 )
);
defparam \top/processor/sha_core/n3629_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [8]),
	.I3(\top/processor/sha_core/w[9] [8]),
	.F(\top/processor/sha_core/n3630_174 )
);
defparam \top/processor/sha_core/n3630_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [7]),
	.I3(\top/processor/sha_core/w[9] [7]),
	.F(\top/processor/sha_core/n3631_174 )
);
defparam \top/processor/sha_core/n3631_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [6]),
	.I3(\top/processor/sha_core/w[9] [6]),
	.F(\top/processor/sha_core/n3632_174 )
);
defparam \top/processor/sha_core/n3632_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [5]),
	.I3(\top/processor/sha_core/w[9] [5]),
	.F(\top/processor/sha_core/n3633_174 )
);
defparam \top/processor/sha_core/n3633_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [4]),
	.I3(\top/processor/sha_core/w[9] [4]),
	.F(\top/processor/sha_core/n3634_174 )
);
defparam \top/processor/sha_core/n3634_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [3]),
	.I3(\top/processor/sha_core/w[9] [3]),
	.F(\top/processor/sha_core/n3635_174 )
);
defparam \top/processor/sha_core/n3635_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [2]),
	.I3(\top/processor/sha_core/w[9] [2]),
	.F(\top/processor/sha_core/n3636_174 )
);
defparam \top/processor/sha_core/n3636_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [1]),
	.I3(\top/processor/sha_core/w[9] [1]),
	.F(\top/processor/sha_core/n3637_174 )
);
defparam \top/processor/sha_core/n3637_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s153  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[11] [0]),
	.I3(\top/processor/sha_core/w[9] [0]),
	.F(\top/processor/sha_core/n3638_174 )
);
defparam \top/processor/sha_core/n3638_s153 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3492_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_119 ),
	.I3(\top/processor/sha_core/n3492_173 ),
	.F(\top/processor/sha_core/n3492_151 )
);
defparam \top/processor/sha_core/n3492_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [27]),
	.I2(\top/processor/sha_core/w[9] [27]),
	.F(\top/processor/sha_core/n3492_152 )
);
defparam \top/processor/sha_core/n3492_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [27]),
	.I2(\top/processor/sha_core/w[13] [27]),
	.F(\top/processor/sha_core/n3492_153 )
);
defparam \top/processor/sha_core/n3492_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_173 ),
	.I3(\top/processor/sha_core/n3492_152 ),
	.F(\top/processor/sha_core/n3864_118 )
);
defparam \top/processor/sha_core/n3864_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [27]),
	.I2(\top/processor/sha_core/w[15] [27]),
	.F(\top/processor/sha_core/n3864_119 )
);
defparam \top/processor/sha_core/n3864_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3492_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_121 ),
	.I3(\top/processor/sha_core/n3492_174 ),
	.F(\top/processor/sha_core/n3492_154 )
);
defparam \top/processor/sha_core/n3492_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [27]),
	.I2(\top/processor/sha_core/w[17] [27]),
	.F(\top/processor/sha_core/n3492_155 )
);
defparam \top/processor/sha_core/n3492_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [27]),
	.I2(\top/processor/sha_core/w[21] [27]),
	.F(\top/processor/sha_core/n3492_156 )
);
defparam \top/processor/sha_core/n3492_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_174 ),
	.I3(\top/processor/sha_core/n3492_155 ),
	.F(\top/processor/sha_core/n3864_120 )
);
defparam \top/processor/sha_core/n3864_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [27]),
	.I2(\top/processor/sha_core/w[23] [27]),
	.F(\top/processor/sha_core/n3864_121 )
);
defparam \top/processor/sha_core/n3864_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [31]),
	.I3(\top/processor/sha_core/w[13] [31]),
	.F(\top/processor/sha_core/n3607_175 )
);
defparam \top/processor/sha_core/n3607_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [30]),
	.I3(\top/processor/sha_core/w[13] [30]),
	.F(\top/processor/sha_core/n3608_175 )
);
defparam \top/processor/sha_core/n3608_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [29]),
	.I3(\top/processor/sha_core/w[13] [29]),
	.F(\top/processor/sha_core/n3609_175 )
);
defparam \top/processor/sha_core/n3609_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [28]),
	.I3(\top/processor/sha_core/w[13] [28]),
	.F(\top/processor/sha_core/n3610_175 )
);
defparam \top/processor/sha_core/n3610_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [27]),
	.I3(\top/processor/sha_core/w[13] [27]),
	.F(\top/processor/sha_core/n3611_175 )
);
defparam \top/processor/sha_core/n3611_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [26]),
	.I3(\top/processor/sha_core/w[13] [26]),
	.F(\top/processor/sha_core/n3612_175 )
);
defparam \top/processor/sha_core/n3612_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [25]),
	.I3(\top/processor/sha_core/w[13] [25]),
	.F(\top/processor/sha_core/n3613_175 )
);
defparam \top/processor/sha_core/n3613_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [24]),
	.I3(\top/processor/sha_core/w[13] [24]),
	.F(\top/processor/sha_core/n3614_175 )
);
defparam \top/processor/sha_core/n3614_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [23]),
	.I3(\top/processor/sha_core/w[13] [23]),
	.F(\top/processor/sha_core/n3615_175 )
);
defparam \top/processor/sha_core/n3615_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [22]),
	.I3(\top/processor/sha_core/w[13] [22]),
	.F(\top/processor/sha_core/n3616_175 )
);
defparam \top/processor/sha_core/n3616_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [21]),
	.I3(\top/processor/sha_core/w[13] [21]),
	.F(\top/processor/sha_core/n3617_175 )
);
defparam \top/processor/sha_core/n3617_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [20]),
	.I3(\top/processor/sha_core/w[13] [20]),
	.F(\top/processor/sha_core/n3618_175 )
);
defparam \top/processor/sha_core/n3618_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [19]),
	.I3(\top/processor/sha_core/w[13] [19]),
	.F(\top/processor/sha_core/n3619_175 )
);
defparam \top/processor/sha_core/n3619_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [18]),
	.I3(\top/processor/sha_core/w[13] [18]),
	.F(\top/processor/sha_core/n3620_175 )
);
defparam \top/processor/sha_core/n3620_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [17]),
	.I3(\top/processor/sha_core/w[13] [17]),
	.F(\top/processor/sha_core/n3621_175 )
);
defparam \top/processor/sha_core/n3621_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3492_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_123 ),
	.I3(\top/processor/sha_core/n3492_175 ),
	.F(\top/processor/sha_core/n3492_157 )
);
defparam \top/processor/sha_core/n3492_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [27]),
	.I2(\top/processor/sha_core/w[25] [27]),
	.F(\top/processor/sha_core/n3492_158 )
);
defparam \top/processor/sha_core/n3492_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [27]),
	.I2(\top/processor/sha_core/w[29] [27]),
	.F(\top/processor/sha_core/n3492_159 )
);
defparam \top/processor/sha_core/n3492_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_175 ),
	.I3(\top/processor/sha_core/n3492_158 ),
	.F(\top/processor/sha_core/n3864_122 )
);
defparam \top/processor/sha_core/n3864_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [27]),
	.I2(\top/processor/sha_core/w[31] [27]),
	.F(\top/processor/sha_core/n3864_123 )
);
defparam \top/processor/sha_core/n3864_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3622_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [16]),
	.I3(\top/processor/sha_core/w[13] [16]),
	.F(\top/processor/sha_core/n3622_175 )
);
defparam \top/processor/sha_core/n3622_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [15]),
	.I3(\top/processor/sha_core/w[13] [15]),
	.F(\top/processor/sha_core/n3623_175 )
);
defparam \top/processor/sha_core/n3623_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [14]),
	.I3(\top/processor/sha_core/w[13] [14]),
	.F(\top/processor/sha_core/n3624_175 )
);
defparam \top/processor/sha_core/n3624_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [13]),
	.I3(\top/processor/sha_core/w[13] [13]),
	.F(\top/processor/sha_core/n3625_175 )
);
defparam \top/processor/sha_core/n3625_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [12]),
	.I3(\top/processor/sha_core/w[13] [12]),
	.F(\top/processor/sha_core/n3626_175 )
);
defparam \top/processor/sha_core/n3626_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [11]),
	.I3(\top/processor/sha_core/w[13] [11]),
	.F(\top/processor/sha_core/n3627_175 )
);
defparam \top/processor/sha_core/n3627_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [10]),
	.I3(\top/processor/sha_core/w[13] [10]),
	.F(\top/processor/sha_core/n3628_175 )
);
defparam \top/processor/sha_core/n3628_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [9]),
	.I3(\top/processor/sha_core/w[13] [9]),
	.F(\top/processor/sha_core/n3629_175 )
);
defparam \top/processor/sha_core/n3629_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [8]),
	.I3(\top/processor/sha_core/w[13] [8]),
	.F(\top/processor/sha_core/n3630_175 )
);
defparam \top/processor/sha_core/n3630_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [7]),
	.I3(\top/processor/sha_core/w[13] [7]),
	.F(\top/processor/sha_core/n3631_175 )
);
defparam \top/processor/sha_core/n3631_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [6]),
	.I3(\top/processor/sha_core/w[13] [6]),
	.F(\top/processor/sha_core/n3632_175 )
);
defparam \top/processor/sha_core/n3632_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [5]),
	.I3(\top/processor/sha_core/w[13] [5]),
	.F(\top/processor/sha_core/n3633_175 )
);
defparam \top/processor/sha_core/n3633_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [4]),
	.I3(\top/processor/sha_core/w[13] [4]),
	.F(\top/processor/sha_core/n3634_175 )
);
defparam \top/processor/sha_core/n3634_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [3]),
	.I3(\top/processor/sha_core/w[13] [3]),
	.F(\top/processor/sha_core/n3635_175 )
);
defparam \top/processor/sha_core/n3635_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [2]),
	.I3(\top/processor/sha_core/w[13] [2]),
	.F(\top/processor/sha_core/n3636_175 )
);
defparam \top/processor/sha_core/n3636_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [1]),
	.I3(\top/processor/sha_core/w[13] [1]),
	.F(\top/processor/sha_core/n3637_175 )
);
defparam \top/processor/sha_core/n3637_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[15] [0]),
	.I3(\top/processor/sha_core/w[13] [0]),
	.F(\top/processor/sha_core/n3638_175 )
);
defparam \top/processor/sha_core/n3638_s154 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3492_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_125 ),
	.I3(\top/processor/sha_core/n3492_176 ),
	.F(\top/processor/sha_core/n3492_160 )
);
defparam \top/processor/sha_core/n3492_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [27]),
	.I2(\top/processor/sha_core/w[33] [27]),
	.F(\top/processor/sha_core/n3492_161 )
);
defparam \top/processor/sha_core/n3492_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [27]),
	.I2(\top/processor/sha_core/w[37] [27]),
	.F(\top/processor/sha_core/n3492_162 )
);
defparam \top/processor/sha_core/n3492_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_176 ),
	.I3(\top/processor/sha_core/n3492_161 ),
	.F(\top/processor/sha_core/n3864_124 )
);
defparam \top/processor/sha_core/n3864_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [27]),
	.I2(\top/processor/sha_core/w[39] [27]),
	.F(\top/processor/sha_core/n3864_125 )
);
defparam \top/processor/sha_core/n3864_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3492_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_127 ),
	.I3(\top/processor/sha_core/n3492_177 ),
	.F(\top/processor/sha_core/n3492_163 )
);
defparam \top/processor/sha_core/n3492_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [27]),
	.I2(\top/processor/sha_core/w[41] [27]),
	.F(\top/processor/sha_core/n3492_164 )
);
defparam \top/processor/sha_core/n3492_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [27]),
	.I2(\top/processor/sha_core/w[45] [27]),
	.F(\top/processor/sha_core/n3492_165 )
);
defparam \top/processor/sha_core/n3492_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_177 ),
	.I3(\top/processor/sha_core/n3492_164 ),
	.F(\top/processor/sha_core/n3864_126 )
);
defparam \top/processor/sha_core/n3864_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [27]),
	.I2(\top/processor/sha_core/w[47] [27]),
	.F(\top/processor/sha_core/n3864_127 )
);
defparam \top/processor/sha_core/n3864_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [31]),
	.I3(\top/processor/sha_core/w[17] [31]),
	.F(\top/processor/sha_core/n3607_176 )
);
defparam \top/processor/sha_core/n3607_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [30]),
	.I3(\top/processor/sha_core/w[17] [30]),
	.F(\top/processor/sha_core/n3608_176 )
);
defparam \top/processor/sha_core/n3608_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [29]),
	.I3(\top/processor/sha_core/w[17] [29]),
	.F(\top/processor/sha_core/n3609_176 )
);
defparam \top/processor/sha_core/n3609_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [28]),
	.I3(\top/processor/sha_core/w[17] [28]),
	.F(\top/processor/sha_core/n3610_176 )
);
defparam \top/processor/sha_core/n3610_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [27]),
	.I3(\top/processor/sha_core/w[17] [27]),
	.F(\top/processor/sha_core/n3611_176 )
);
defparam \top/processor/sha_core/n3611_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [26]),
	.I3(\top/processor/sha_core/w[17] [26]),
	.F(\top/processor/sha_core/n3612_176 )
);
defparam \top/processor/sha_core/n3612_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [25]),
	.I3(\top/processor/sha_core/w[17] [25]),
	.F(\top/processor/sha_core/n3613_176 )
);
defparam \top/processor/sha_core/n3613_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [24]),
	.I3(\top/processor/sha_core/w[17] [24]),
	.F(\top/processor/sha_core/n3614_176 )
);
defparam \top/processor/sha_core/n3614_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [23]),
	.I3(\top/processor/sha_core/w[17] [23]),
	.F(\top/processor/sha_core/n3615_176 )
);
defparam \top/processor/sha_core/n3615_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [22]),
	.I3(\top/processor/sha_core/w[17] [22]),
	.F(\top/processor/sha_core/n3616_176 )
);
defparam \top/processor/sha_core/n3616_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [21]),
	.I3(\top/processor/sha_core/w[17] [21]),
	.F(\top/processor/sha_core/n3617_176 )
);
defparam \top/processor/sha_core/n3617_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3492_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_129 ),
	.I3(\top/processor/sha_core/n3492_178 ),
	.F(\top/processor/sha_core/n3492_166 )
);
defparam \top/processor/sha_core/n3492_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [27]),
	.I2(\top/processor/sha_core/w[49] [27]),
	.F(\top/processor/sha_core/n3492_167 )
);
defparam \top/processor/sha_core/n3492_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [27]),
	.I2(\top/processor/sha_core/w[53] [27]),
	.F(\top/processor/sha_core/n3492_168 )
);
defparam \top/processor/sha_core/n3492_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_178 ),
	.I3(\top/processor/sha_core/n3492_167 ),
	.F(\top/processor/sha_core/n3864_128 )
);
defparam \top/processor/sha_core/n3864_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [27]),
	.I2(\top/processor/sha_core/w[55] [27]),
	.F(\top/processor/sha_core/n3864_129 )
);
defparam \top/processor/sha_core/n3864_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3618_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [20]),
	.I3(\top/processor/sha_core/w[17] [20]),
	.F(\top/processor/sha_core/n3618_176 )
);
defparam \top/processor/sha_core/n3618_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [19]),
	.I3(\top/processor/sha_core/w[17] [19]),
	.F(\top/processor/sha_core/n3619_176 )
);
defparam \top/processor/sha_core/n3619_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [18]),
	.I3(\top/processor/sha_core/w[17] [18]),
	.F(\top/processor/sha_core/n3620_176 )
);
defparam \top/processor/sha_core/n3620_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [17]),
	.I3(\top/processor/sha_core/w[17] [17]),
	.F(\top/processor/sha_core/n3621_176 )
);
defparam \top/processor/sha_core/n3621_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [16]),
	.I3(\top/processor/sha_core/w[17] [16]),
	.F(\top/processor/sha_core/n3622_176 )
);
defparam \top/processor/sha_core/n3622_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [15]),
	.I3(\top/processor/sha_core/w[17] [15]),
	.F(\top/processor/sha_core/n3623_176 )
);
defparam \top/processor/sha_core/n3623_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [14]),
	.I3(\top/processor/sha_core/w[17] [14]),
	.F(\top/processor/sha_core/n3624_176 )
);
defparam \top/processor/sha_core/n3624_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [13]),
	.I3(\top/processor/sha_core/w[17] [13]),
	.F(\top/processor/sha_core/n3625_176 )
);
defparam \top/processor/sha_core/n3625_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [12]),
	.I3(\top/processor/sha_core/w[17] [12]),
	.F(\top/processor/sha_core/n3626_176 )
);
defparam \top/processor/sha_core/n3626_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [11]),
	.I3(\top/processor/sha_core/w[17] [11]),
	.F(\top/processor/sha_core/n3627_176 )
);
defparam \top/processor/sha_core/n3627_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [10]),
	.I3(\top/processor/sha_core/w[17] [10]),
	.F(\top/processor/sha_core/n3628_176 )
);
defparam \top/processor/sha_core/n3628_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [9]),
	.I3(\top/processor/sha_core/w[17] [9]),
	.F(\top/processor/sha_core/n3629_176 )
);
defparam \top/processor/sha_core/n3629_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [8]),
	.I3(\top/processor/sha_core/w[17] [8]),
	.F(\top/processor/sha_core/n3630_176 )
);
defparam \top/processor/sha_core/n3630_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [7]),
	.I3(\top/processor/sha_core/w[17] [7]),
	.F(\top/processor/sha_core/n3631_176 )
);
defparam \top/processor/sha_core/n3631_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [6]),
	.I3(\top/processor/sha_core/w[17] [6]),
	.F(\top/processor/sha_core/n3632_176 )
);
defparam \top/processor/sha_core/n3632_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [5]),
	.I3(\top/processor/sha_core/w[17] [5]),
	.F(\top/processor/sha_core/n3633_176 )
);
defparam \top/processor/sha_core/n3633_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [4]),
	.I3(\top/processor/sha_core/w[17] [4]),
	.F(\top/processor/sha_core/n3634_176 )
);
defparam \top/processor/sha_core/n3634_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [3]),
	.I3(\top/processor/sha_core/w[17] [3]),
	.F(\top/processor/sha_core/n3635_176 )
);
defparam \top/processor/sha_core/n3635_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [2]),
	.I3(\top/processor/sha_core/w[17] [2]),
	.F(\top/processor/sha_core/n3636_176 )
);
defparam \top/processor/sha_core/n3636_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [1]),
	.I3(\top/processor/sha_core/w[17] [1]),
	.F(\top/processor/sha_core/n3637_176 )
);
defparam \top/processor/sha_core/n3637_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3492_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3864_131 ),
	.I3(\top/processor/sha_core/n3492_179 ),
	.F(\top/processor/sha_core/n3492_169 )
);
defparam \top/processor/sha_core/n3492_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3492_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [27]),
	.I2(\top/processor/sha_core/w[57] [27]),
	.F(\top/processor/sha_core/n3492_170 )
);
defparam \top/processor/sha_core/n3492_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [27]),
	.I2(\top/processor/sha_core/w[61] [27]),
	.F(\top/processor/sha_core/n3492_171 )
);
defparam \top/processor/sha_core/n3492_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3864_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3492_179 ),
	.I3(\top/processor/sha_core/n3492_170 ),
	.F(\top/processor/sha_core/n3864_130 )
);
defparam \top/processor/sha_core/n3864_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3864_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [27]),
	.I2(\top/processor/sha_core/w[63] [27]),
	.F(\top/processor/sha_core/n3864_131 )
);
defparam \top/processor/sha_core/n3864_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_129 ),
	.I3(\top/processor/sha_core/n3488_178 ),
	.F(\top/processor/sha_core/n3488_166 )
);
defparam \top/processor/sha_core/n3488_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [31]),
	.I2(\top/processor/sha_core/w[25] [31]),
	.F(\top/processor/sha_core/n3488_167 )
);
defparam \top/processor/sha_core/n3488_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [31]),
	.I2(\top/processor/sha_core/w[29] [31]),
	.F(\top/processor/sha_core/n3488_168 )
);
defparam \top/processor/sha_core/n3488_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_178 ),
	.I3(\top/processor/sha_core/n3488_167 ),
	.F(\top/processor/sha_core/n3860_128 )
);
defparam \top/processor/sha_core/n3860_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3860_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [31]),
	.I2(\top/processor/sha_core/w[31] [31]),
	.F(\top/processor/sha_core/n3860_129 )
);
defparam \top/processor/sha_core/n3860_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3638_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[19] [0]),
	.I3(\top/processor/sha_core/w[17] [0]),
	.F(\top/processor/sha_core/n3638_176 )
);
defparam \top/processor/sha_core/n3638_s155 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s135  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_117 ),
	.I3(\top/processor/sha_core/n3493_172 ),
	.F(\top/processor/sha_core/n3493_148 )
);
defparam \top/processor/sha_core/n3493_s135 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s136  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [26]),
	.I2(\top/processor/sha_core/w[1] [26]),
	.F(\top/processor/sha_core/n3493_149 )
);
defparam \top/processor/sha_core/n3493_s136 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s137  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [26]),
	.I2(\top/processor/sha_core/w[5] [26]),
	.F(\top/processor/sha_core/n3493_150 )
);
defparam \top/processor/sha_core/n3493_s137 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s103  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_172 ),
	.I3(\top/processor/sha_core/n3493_149 ),
	.F(\top/processor/sha_core/n3865_116 )
);
defparam \top/processor/sha_core/n3865_s103 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s104  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [26]),
	.I2(\top/processor/sha_core/w[7] [26]),
	.F(\top/processor/sha_core/n3865_117 )
);
defparam \top/processor/sha_core/n3865_s104 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [31]),
	.I3(\top/processor/sha_core/w[21] [31]),
	.F(\top/processor/sha_core/n3607_177 )
);
defparam \top/processor/sha_core/n3607_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [30]),
	.I3(\top/processor/sha_core/w[21] [30]),
	.F(\top/processor/sha_core/n3608_177 )
);
defparam \top/processor/sha_core/n3608_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [29]),
	.I3(\top/processor/sha_core/w[21] [29]),
	.F(\top/processor/sha_core/n3609_177 )
);
defparam \top/processor/sha_core/n3609_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [28]),
	.I3(\top/processor/sha_core/w[21] [28]),
	.F(\top/processor/sha_core/n3610_177 )
);
defparam \top/processor/sha_core/n3610_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [27]),
	.I3(\top/processor/sha_core/w[21] [27]),
	.F(\top/processor/sha_core/n3611_177 )
);
defparam \top/processor/sha_core/n3611_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [26]),
	.I3(\top/processor/sha_core/w[21] [26]),
	.F(\top/processor/sha_core/n3612_177 )
);
defparam \top/processor/sha_core/n3612_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [25]),
	.I3(\top/processor/sha_core/w[21] [25]),
	.F(\top/processor/sha_core/n3613_177 )
);
defparam \top/processor/sha_core/n3613_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s138  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_119 ),
	.I3(\top/processor/sha_core/n3493_173 ),
	.F(\top/processor/sha_core/n3493_151 )
);
defparam \top/processor/sha_core/n3493_s138 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s139  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [26]),
	.I2(\top/processor/sha_core/w[9] [26]),
	.F(\top/processor/sha_core/n3493_152 )
);
defparam \top/processor/sha_core/n3493_s139 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s140  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [26]),
	.I2(\top/processor/sha_core/w[13] [26]),
	.F(\top/processor/sha_core/n3493_153 )
);
defparam \top/processor/sha_core/n3493_s140 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s105  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_173 ),
	.I3(\top/processor/sha_core/n3493_152 ),
	.F(\top/processor/sha_core/n3865_118 )
);
defparam \top/processor/sha_core/n3865_s105 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s106  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [26]),
	.I2(\top/processor/sha_core/w[15] [26]),
	.F(\top/processor/sha_core/n3865_119 )
);
defparam \top/processor/sha_core/n3865_s106 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3614_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [24]),
	.I3(\top/processor/sha_core/w[21] [24]),
	.F(\top/processor/sha_core/n3614_177 )
);
defparam \top/processor/sha_core/n3614_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [23]),
	.I3(\top/processor/sha_core/w[21] [23]),
	.F(\top/processor/sha_core/n3615_177 )
);
defparam \top/processor/sha_core/n3615_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [22]),
	.I3(\top/processor/sha_core/w[21] [22]),
	.F(\top/processor/sha_core/n3616_177 )
);
defparam \top/processor/sha_core/n3616_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [21]),
	.I3(\top/processor/sha_core/w[21] [21]),
	.F(\top/processor/sha_core/n3617_177 )
);
defparam \top/processor/sha_core/n3617_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [20]),
	.I3(\top/processor/sha_core/w[21] [20]),
	.F(\top/processor/sha_core/n3618_177 )
);
defparam \top/processor/sha_core/n3618_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [19]),
	.I3(\top/processor/sha_core/w[21] [19]),
	.F(\top/processor/sha_core/n3619_177 )
);
defparam \top/processor/sha_core/n3619_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [18]),
	.I3(\top/processor/sha_core/w[21] [18]),
	.F(\top/processor/sha_core/n3620_177 )
);
defparam \top/processor/sha_core/n3620_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [17]),
	.I3(\top/processor/sha_core/w[21] [17]),
	.F(\top/processor/sha_core/n3621_177 )
);
defparam \top/processor/sha_core/n3621_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [16]),
	.I3(\top/processor/sha_core/w[21] [16]),
	.F(\top/processor/sha_core/n3622_177 )
);
defparam \top/processor/sha_core/n3622_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [15]),
	.I3(\top/processor/sha_core/w[21] [15]),
	.F(\top/processor/sha_core/n3623_177 )
);
defparam \top/processor/sha_core/n3623_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [14]),
	.I3(\top/processor/sha_core/w[21] [14]),
	.F(\top/processor/sha_core/n3624_177 )
);
defparam \top/processor/sha_core/n3624_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [13]),
	.I3(\top/processor/sha_core/w[21] [13]),
	.F(\top/processor/sha_core/n3625_177 )
);
defparam \top/processor/sha_core/n3625_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [12]),
	.I3(\top/processor/sha_core/w[21] [12]),
	.F(\top/processor/sha_core/n3626_177 )
);
defparam \top/processor/sha_core/n3626_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [11]),
	.I3(\top/processor/sha_core/w[21] [11]),
	.F(\top/processor/sha_core/n3627_177 )
);
defparam \top/processor/sha_core/n3627_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [10]),
	.I3(\top/processor/sha_core/w[21] [10]),
	.F(\top/processor/sha_core/n3628_177 )
);
defparam \top/processor/sha_core/n3628_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [9]),
	.I3(\top/processor/sha_core/w[21] [9]),
	.F(\top/processor/sha_core/n3629_177 )
);
defparam \top/processor/sha_core/n3629_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [8]),
	.I3(\top/processor/sha_core/w[21] [8]),
	.F(\top/processor/sha_core/n3630_177 )
);
defparam \top/processor/sha_core/n3630_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [7]),
	.I3(\top/processor/sha_core/w[21] [7]),
	.F(\top/processor/sha_core/n3631_177 )
);
defparam \top/processor/sha_core/n3631_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [6]),
	.I3(\top/processor/sha_core/w[21] [6]),
	.F(\top/processor/sha_core/n3632_177 )
);
defparam \top/processor/sha_core/n3632_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [5]),
	.I3(\top/processor/sha_core/w[21] [5]),
	.F(\top/processor/sha_core/n3633_177 )
);
defparam \top/processor/sha_core/n3633_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s141  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_121 ),
	.I3(\top/processor/sha_core/n3493_174 ),
	.F(\top/processor/sha_core/n3493_154 )
);
defparam \top/processor/sha_core/n3493_s141 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s142  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[16] [26]),
	.I2(\top/processor/sha_core/w[17] [26]),
	.F(\top/processor/sha_core/n3493_155 )
);
defparam \top/processor/sha_core/n3493_s142 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s143  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[20] [26]),
	.I2(\top/processor/sha_core/w[21] [26]),
	.F(\top/processor/sha_core/n3493_156 )
);
defparam \top/processor/sha_core/n3493_s143 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s107  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_174 ),
	.I3(\top/processor/sha_core/n3493_155 ),
	.F(\top/processor/sha_core/n3865_120 )
);
defparam \top/processor/sha_core/n3865_s107 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s108  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[22] [26]),
	.I2(\top/processor/sha_core/w[23] [26]),
	.F(\top/processor/sha_core/n3865_121 )
);
defparam \top/processor/sha_core/n3865_s108 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3634_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [4]),
	.I3(\top/processor/sha_core/w[21] [4]),
	.F(\top/processor/sha_core/n3634_177 )
);
defparam \top/processor/sha_core/n3634_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [3]),
	.I3(\top/processor/sha_core/w[21] [3]),
	.F(\top/processor/sha_core/n3635_177 )
);
defparam \top/processor/sha_core/n3635_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [2]),
	.I3(\top/processor/sha_core/w[21] [2]),
	.F(\top/processor/sha_core/n3636_177 )
);
defparam \top/processor/sha_core/n3636_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [1]),
	.I3(\top/processor/sha_core/w[21] [1]),
	.F(\top/processor/sha_core/n3637_177 )
);
defparam \top/processor/sha_core/n3637_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s156  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[23] [0]),
	.I3(\top/processor/sha_core/w[21] [0]),
	.F(\top/processor/sha_core/n3638_177 )
);
defparam \top/processor/sha_core/n3638_s156 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s144  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_123 ),
	.I3(\top/processor/sha_core/n3493_175 ),
	.F(\top/processor/sha_core/n3493_157 )
);
defparam \top/processor/sha_core/n3493_s144 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s145  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[24] [26]),
	.I2(\top/processor/sha_core/w[25] [26]),
	.F(\top/processor/sha_core/n3493_158 )
);
defparam \top/processor/sha_core/n3493_s145 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s146  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[28] [26]),
	.I2(\top/processor/sha_core/w[29] [26]),
	.F(\top/processor/sha_core/n3493_159 )
);
defparam \top/processor/sha_core/n3493_s146 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s109  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_175 ),
	.I3(\top/processor/sha_core/n3493_158 ),
	.F(\top/processor/sha_core/n3865_122 )
);
defparam \top/processor/sha_core/n3865_s109 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s110  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[30] [26]),
	.I2(\top/processor/sha_core/w[31] [26]),
	.F(\top/processor/sha_core/n3865_123 )
);
defparam \top/processor/sha_core/n3865_s110 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [31]),
	.I3(\top/processor/sha_core/w[25] [31]),
	.F(\top/processor/sha_core/n3607_178 )
);
defparam \top/processor/sha_core/n3607_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [30]),
	.I3(\top/processor/sha_core/w[25] [30]),
	.F(\top/processor/sha_core/n3608_178 )
);
defparam \top/processor/sha_core/n3608_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [29]),
	.I3(\top/processor/sha_core/w[25] [29]),
	.F(\top/processor/sha_core/n3609_178 )
);
defparam \top/processor/sha_core/n3609_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s147  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_125 ),
	.I3(\top/processor/sha_core/n3493_176 ),
	.F(\top/processor/sha_core/n3493_160 )
);
defparam \top/processor/sha_core/n3493_s147 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s148  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [26]),
	.I2(\top/processor/sha_core/w[33] [26]),
	.F(\top/processor/sha_core/n3493_161 )
);
defparam \top/processor/sha_core/n3493_s148 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s149  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [26]),
	.I2(\top/processor/sha_core/w[37] [26]),
	.F(\top/processor/sha_core/n3493_162 )
);
defparam \top/processor/sha_core/n3493_s149 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s111  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_176 ),
	.I3(\top/processor/sha_core/n3493_161 ),
	.F(\top/processor/sha_core/n3865_124 )
);
defparam \top/processor/sha_core/n3865_s111 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s112  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [26]),
	.I2(\top/processor/sha_core/w[39] [26]),
	.F(\top/processor/sha_core/n3865_125 )
);
defparam \top/processor/sha_core/n3865_s112 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3610_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [28]),
	.I3(\top/processor/sha_core/w[25] [28]),
	.F(\top/processor/sha_core/n3610_178 )
);
defparam \top/processor/sha_core/n3610_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [27]),
	.I3(\top/processor/sha_core/w[25] [27]),
	.F(\top/processor/sha_core/n3611_178 )
);
defparam \top/processor/sha_core/n3611_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [26]),
	.I3(\top/processor/sha_core/w[25] [26]),
	.F(\top/processor/sha_core/n3612_178 )
);
defparam \top/processor/sha_core/n3612_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [25]),
	.I3(\top/processor/sha_core/w[25] [25]),
	.F(\top/processor/sha_core/n3613_178 )
);
defparam \top/processor/sha_core/n3613_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [24]),
	.I3(\top/processor/sha_core/w[25] [24]),
	.F(\top/processor/sha_core/n3614_178 )
);
defparam \top/processor/sha_core/n3614_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [23]),
	.I3(\top/processor/sha_core/w[25] [23]),
	.F(\top/processor/sha_core/n3615_178 )
);
defparam \top/processor/sha_core/n3615_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [22]),
	.I3(\top/processor/sha_core/w[25] [22]),
	.F(\top/processor/sha_core/n3616_178 )
);
defparam \top/processor/sha_core/n3616_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [21]),
	.I3(\top/processor/sha_core/w[25] [21]),
	.F(\top/processor/sha_core/n3617_178 )
);
defparam \top/processor/sha_core/n3617_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [20]),
	.I3(\top/processor/sha_core/w[25] [20]),
	.F(\top/processor/sha_core/n3618_178 )
);
defparam \top/processor/sha_core/n3618_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [19]),
	.I3(\top/processor/sha_core/w[25] [19]),
	.F(\top/processor/sha_core/n3619_178 )
);
defparam \top/processor/sha_core/n3619_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [18]),
	.I3(\top/processor/sha_core/w[25] [18]),
	.F(\top/processor/sha_core/n3620_178 )
);
defparam \top/processor/sha_core/n3620_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [17]),
	.I3(\top/processor/sha_core/w[25] [17]),
	.F(\top/processor/sha_core/n3621_178 )
);
defparam \top/processor/sha_core/n3621_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [16]),
	.I3(\top/processor/sha_core/w[25] [16]),
	.F(\top/processor/sha_core/n3622_178 )
);
defparam \top/processor/sha_core/n3622_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [15]),
	.I3(\top/processor/sha_core/w[25] [15]),
	.F(\top/processor/sha_core/n3623_178 )
);
defparam \top/processor/sha_core/n3623_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [14]),
	.I3(\top/processor/sha_core/w[25] [14]),
	.F(\top/processor/sha_core/n3624_178 )
);
defparam \top/processor/sha_core/n3624_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [13]),
	.I3(\top/processor/sha_core/w[25] [13]),
	.F(\top/processor/sha_core/n3625_178 )
);
defparam \top/processor/sha_core/n3625_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3626_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [12]),
	.I3(\top/processor/sha_core/w[25] [12]),
	.F(\top/processor/sha_core/n3626_178 )
);
defparam \top/processor/sha_core/n3626_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [11]),
	.I3(\top/processor/sha_core/w[25] [11]),
	.F(\top/processor/sha_core/n3627_178 )
);
defparam \top/processor/sha_core/n3627_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [10]),
	.I3(\top/processor/sha_core/w[25] [10]),
	.F(\top/processor/sha_core/n3628_178 )
);
defparam \top/processor/sha_core/n3628_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [9]),
	.I3(\top/processor/sha_core/w[25] [9]),
	.F(\top/processor/sha_core/n3629_178 )
);
defparam \top/processor/sha_core/n3629_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s150  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_127 ),
	.I3(\top/processor/sha_core/n3493_177 ),
	.F(\top/processor/sha_core/n3493_163 )
);
defparam \top/processor/sha_core/n3493_s150 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s151  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[40] [26]),
	.I2(\top/processor/sha_core/w[41] [26]),
	.F(\top/processor/sha_core/n3493_164 )
);
defparam \top/processor/sha_core/n3493_s151 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s152  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[44] [26]),
	.I2(\top/processor/sha_core/w[45] [26]),
	.F(\top/processor/sha_core/n3493_165 )
);
defparam \top/processor/sha_core/n3493_s152 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s113  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_177 ),
	.I3(\top/processor/sha_core/n3493_164 ),
	.F(\top/processor/sha_core/n3865_126 )
);
defparam \top/processor/sha_core/n3865_s113 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s114  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[46] [26]),
	.I2(\top/processor/sha_core/w[47] [26]),
	.F(\top/processor/sha_core/n3865_127 )
);
defparam \top/processor/sha_core/n3865_s114 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3630_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [8]),
	.I3(\top/processor/sha_core/w[25] [8]),
	.F(\top/processor/sha_core/n3630_178 )
);
defparam \top/processor/sha_core/n3630_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [7]),
	.I3(\top/processor/sha_core/w[25] [7]),
	.F(\top/processor/sha_core/n3631_178 )
);
defparam \top/processor/sha_core/n3631_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [6]),
	.I3(\top/processor/sha_core/w[25] [6]),
	.F(\top/processor/sha_core/n3632_178 )
);
defparam \top/processor/sha_core/n3632_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [5]),
	.I3(\top/processor/sha_core/w[25] [5]),
	.F(\top/processor/sha_core/n3633_178 )
);
defparam \top/processor/sha_core/n3633_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [4]),
	.I3(\top/processor/sha_core/w[25] [4]),
	.F(\top/processor/sha_core/n3634_178 )
);
defparam \top/processor/sha_core/n3634_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [3]),
	.I3(\top/processor/sha_core/w[25] [3]),
	.F(\top/processor/sha_core/n3635_178 )
);
defparam \top/processor/sha_core/n3635_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [2]),
	.I3(\top/processor/sha_core/w[25] [2]),
	.F(\top/processor/sha_core/n3636_178 )
);
defparam \top/processor/sha_core/n3636_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [1]),
	.I3(\top/processor/sha_core/w[25] [1]),
	.F(\top/processor/sha_core/n3637_178 )
);
defparam \top/processor/sha_core/n3637_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[27] [0]),
	.I3(\top/processor/sha_core/w[25] [0]),
	.F(\top/processor/sha_core/n3638_178 )
);
defparam \top/processor/sha_core/n3638_s157 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3493_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_129 ),
	.I3(\top/processor/sha_core/n3493_178 ),
	.F(\top/processor/sha_core/n3493_166 )
);
defparam \top/processor/sha_core/n3493_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[48] [26]),
	.I2(\top/processor/sha_core/w[49] [26]),
	.F(\top/processor/sha_core/n3493_167 )
);
defparam \top/processor/sha_core/n3493_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[52] [26]),
	.I2(\top/processor/sha_core/w[53] [26]),
	.F(\top/processor/sha_core/n3493_168 )
);
defparam \top/processor/sha_core/n3493_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_178 ),
	.I3(\top/processor/sha_core/n3493_167 ),
	.F(\top/processor/sha_core/n3865_128 )
);
defparam \top/processor/sha_core/n3865_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[54] [26]),
	.I2(\top/processor/sha_core/w[55] [26]),
	.F(\top/processor/sha_core/n3865_129 )
);
defparam \top/processor/sha_core/n3865_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3493_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3865_131 ),
	.I3(\top/processor/sha_core/n3493_179 ),
	.F(\top/processor/sha_core/n3493_169 )
);
defparam \top/processor/sha_core/n3493_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3493_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[56] [26]),
	.I2(\top/processor/sha_core/w[57] [26]),
	.F(\top/processor/sha_core/n3493_170 )
);
defparam \top/processor/sha_core/n3493_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[60] [26]),
	.I2(\top/processor/sha_core/w[61] [26]),
	.F(\top/processor/sha_core/n3493_171 )
);
defparam \top/processor/sha_core/n3493_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3865_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3493_179 ),
	.I3(\top/processor/sha_core/n3493_170 ),
	.F(\top/processor/sha_core/n3865_130 )
);
defparam \top/processor/sha_core/n3865_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3865_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[62] [26]),
	.I2(\top/processor/sha_core/w[63] [26]),
	.F(\top/processor/sha_core/n3865_131 )
);
defparam \top/processor/sha_core/n3865_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3607_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [31]),
	.I3(\top/processor/sha_core/w[29] [31]),
	.F(\top/processor/sha_core/n3607_179 )
);
defparam \top/processor/sha_core/n3607_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3608_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [30]),
	.I3(\top/processor/sha_core/w[29] [30]),
	.F(\top/processor/sha_core/n3608_179 )
);
defparam \top/processor/sha_core/n3608_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3609_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [29]),
	.I3(\top/processor/sha_core/w[29] [29]),
	.F(\top/processor/sha_core/n3609_179 )
);
defparam \top/processor/sha_core/n3609_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3610_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [28]),
	.I3(\top/processor/sha_core/w[29] [28]),
	.F(\top/processor/sha_core/n3610_179 )
);
defparam \top/processor/sha_core/n3610_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3611_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [27]),
	.I3(\top/processor/sha_core/w[29] [27]),
	.F(\top/processor/sha_core/n3611_179 )
);
defparam \top/processor/sha_core/n3611_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3612_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [26]),
	.I3(\top/processor/sha_core/w[29] [26]),
	.F(\top/processor/sha_core/n3612_179 )
);
defparam \top/processor/sha_core/n3612_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3613_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [25]),
	.I3(\top/processor/sha_core/w[29] [25]),
	.F(\top/processor/sha_core/n3613_179 )
);
defparam \top/processor/sha_core/n3613_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3614_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [24]),
	.I3(\top/processor/sha_core/w[29] [24]),
	.F(\top/processor/sha_core/n3614_179 )
);
defparam \top/processor/sha_core/n3614_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3615_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [23]),
	.I3(\top/processor/sha_core/w[29] [23]),
	.F(\top/processor/sha_core/n3615_179 )
);
defparam \top/processor/sha_core/n3615_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3616_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [22]),
	.I3(\top/processor/sha_core/w[29] [22]),
	.F(\top/processor/sha_core/n3616_179 )
);
defparam \top/processor/sha_core/n3616_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3617_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [21]),
	.I3(\top/processor/sha_core/w[29] [21]),
	.F(\top/processor/sha_core/n3617_179 )
);
defparam \top/processor/sha_core/n3617_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3618_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [20]),
	.I3(\top/processor/sha_core/w[29] [20]),
	.F(\top/processor/sha_core/n3618_179 )
);
defparam \top/processor/sha_core/n3618_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3619_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [19]),
	.I3(\top/processor/sha_core/w[29] [19]),
	.F(\top/processor/sha_core/n3619_179 )
);
defparam \top/processor/sha_core/n3619_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3620_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [18]),
	.I3(\top/processor/sha_core/w[29] [18]),
	.F(\top/processor/sha_core/n3620_179 )
);
defparam \top/processor/sha_core/n3620_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3621_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [17]),
	.I3(\top/processor/sha_core/w[29] [17]),
	.F(\top/processor/sha_core/n3621_179 )
);
defparam \top/processor/sha_core/n3621_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3622_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [16]),
	.I3(\top/processor/sha_core/w[29] [16]),
	.F(\top/processor/sha_core/n3622_179 )
);
defparam \top/processor/sha_core/n3622_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3623_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [15]),
	.I3(\top/processor/sha_core/w[29] [15]),
	.F(\top/processor/sha_core/n3623_179 )
);
defparam \top/processor/sha_core/n3623_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3624_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [14]),
	.I3(\top/processor/sha_core/w[29] [14]),
	.F(\top/processor/sha_core/n3624_179 )
);
defparam \top/processor/sha_core/n3624_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3625_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [13]),
	.I3(\top/processor/sha_core/w[29] [13]),
	.F(\top/processor/sha_core/n3625_179 )
);
defparam \top/processor/sha_core/n3625_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3494_s153  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_129 ),
	.I3(\top/processor/sha_core/n3494_179 ),
	.F(\top/processor/sha_core/n3494_167 )
);
defparam \top/processor/sha_core/n3494_s153 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s154  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[0] [25]),
	.I2(\top/processor/sha_core/w[1] [25]),
	.F(\top/processor/sha_core/n3494_168 )
);
defparam \top/processor/sha_core/n3494_s154 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s155  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[4] [25]),
	.I2(\top/processor/sha_core/w[5] [25]),
	.F(\top/processor/sha_core/n3494_169 )
);
defparam \top/processor/sha_core/n3494_s155 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s115  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_179 ),
	.I3(\top/processor/sha_core/n3494_168 ),
	.F(\top/processor/sha_core/n3866_128 )
);
defparam \top/processor/sha_core/n3866_s115 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s116  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[6] [25]),
	.I2(\top/processor/sha_core/w[7] [25]),
	.F(\top/processor/sha_core/n3866_129 )
);
defparam \top/processor/sha_core/n3866_s116 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3626_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [12]),
	.I3(\top/processor/sha_core/w[29] [12]),
	.F(\top/processor/sha_core/n3626_179 )
);
defparam \top/processor/sha_core/n3626_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3627_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [11]),
	.I3(\top/processor/sha_core/w[29] [11]),
	.F(\top/processor/sha_core/n3627_179 )
);
defparam \top/processor/sha_core/n3627_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3628_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [10]),
	.I3(\top/processor/sha_core/w[29] [10]),
	.F(\top/processor/sha_core/n3628_179 )
);
defparam \top/processor/sha_core/n3628_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3629_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [9]),
	.I3(\top/processor/sha_core/w[29] [9]),
	.F(\top/processor/sha_core/n3629_179 )
);
defparam \top/processor/sha_core/n3629_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3630_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [8]),
	.I3(\top/processor/sha_core/w[29] [8]),
	.F(\top/processor/sha_core/n3630_179 )
);
defparam \top/processor/sha_core/n3630_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3631_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [7]),
	.I3(\top/processor/sha_core/w[29] [7]),
	.F(\top/processor/sha_core/n3631_179 )
);
defparam \top/processor/sha_core/n3631_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3632_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [6]),
	.I3(\top/processor/sha_core/w[29] [6]),
	.F(\top/processor/sha_core/n3632_179 )
);
defparam \top/processor/sha_core/n3632_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3633_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [5]),
	.I3(\top/processor/sha_core/w[29] [5]),
	.F(\top/processor/sha_core/n3633_179 )
);
defparam \top/processor/sha_core/n3633_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3634_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [4]),
	.I3(\top/processor/sha_core/w[29] [4]),
	.F(\top/processor/sha_core/n3634_179 )
);
defparam \top/processor/sha_core/n3634_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3635_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [3]),
	.I3(\top/processor/sha_core/w[29] [3]),
	.F(\top/processor/sha_core/n3635_179 )
);
defparam \top/processor/sha_core/n3635_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3636_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [2]),
	.I3(\top/processor/sha_core/w[29] [2]),
	.F(\top/processor/sha_core/n3636_179 )
);
defparam \top/processor/sha_core/n3636_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3637_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [1]),
	.I3(\top/processor/sha_core/w[29] [1]),
	.F(\top/processor/sha_core/n3637_179 )
);
defparam \top/processor/sha_core/n3637_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3638_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/n3453_7 ),
	.I2(\top/processor/sha_core/w[31] [0]),
	.I3(\top/processor/sha_core/w[29] [0]),
	.F(\top/processor/sha_core/n3638_179 )
);
defparam \top/processor/sha_core/n3638_s158 .INIT=16'h8C9D;
LUT4 \top/processor/sha_core/n3494_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3866_131 ),
	.I3(\top/processor/sha_core/n3494_180 ),
	.F(\top/processor/sha_core/n3494_170 )
);
defparam \top/processor/sha_core/n3494_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3494_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[8] [25]),
	.I2(\top/processor/sha_core/w[9] [25]),
	.F(\top/processor/sha_core/n3494_171 )
);
defparam \top/processor/sha_core/n3494_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[12] [25]),
	.I2(\top/processor/sha_core/w[13] [25]),
	.F(\top/processor/sha_core/n3494_172 )
);
defparam \top/processor/sha_core/n3494_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3866_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3494_180 ),
	.I3(\top/processor/sha_core/n3494_171 ),
	.F(\top/processor/sha_core/n3866_130 )
);
defparam \top/processor/sha_core/n3866_s117 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3866_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[14] [25]),
	.I2(\top/processor/sha_core/w[15] [25]),
	.F(\top/processor/sha_core/n3866_131 )
);
defparam \top/processor/sha_core/n3866_s118 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3488_s156  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/n3462_11 ),
	.I2(\top/processor/sha_core/n3860_131 ),
	.I3(\top/processor/sha_core/n3488_179 ),
	.F(\top/processor/sha_core/n3488_169 )
);
defparam \top/processor/sha_core/n3488_s156 .INIT=16'hD9C8;
LUT3 \top/processor/sha_core/n3488_s157  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[32] [31]),
	.I2(\top/processor/sha_core/w[33] [31]),
	.F(\top/processor/sha_core/n3488_170 )
);
defparam \top/processor/sha_core/n3488_s157 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s158  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[36] [31]),
	.I2(\top/processor/sha_core/w[37] [31]),
	.F(\top/processor/sha_core/n3488_171 )
);
defparam \top/processor/sha_core/n3488_s158 .INIT=8'hE4;
LUT4 \top/processor/sha_core/n3860_s117  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/n3488_179 ),
	.I3(\top/processor/sha_core/n3488_170 ),
	.F(\top/processor/sha_core/n3860_130 )
);
defparam \top/processor/sha_core/n3860_s117 .INIT=16'h8C9D;
LUT3 \top/processor/sha_core/n3860_s118  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[38] [31]),
	.I2(\top/processor/sha_core/w[39] [31]),
	.F(\top/processor/sha_core/n3860_131 )
);
defparam \top/processor/sha_core/n3860_s118 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [25]),
	.I2(\top/processor/sha_core/w[19] [25]),
	.F(\top/processor/sha_core/n3494_173 )
);
defparam \top/processor/sha_core/n3494_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [25]),
	.I2(\top/processor/sha_core/w[27] [25]),
	.F(\top/processor/sha_core/n3494_174 )
);
defparam \top/processor/sha_core/n3494_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [25]),
	.I2(\top/processor/sha_core/w[35] [25]),
	.F(\top/processor/sha_core/n3494_175 )
);
defparam \top/processor/sha_core/n3494_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [25]),
	.I2(\top/processor/sha_core/w[43] [25]),
	.F(\top/processor/sha_core/n3494_176 )
);
defparam \top/processor/sha_core/n3494_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [25]),
	.I2(\top/processor/sha_core/w[51] [25]),
	.F(\top/processor/sha_core/n3494_177 )
);
defparam \top/processor/sha_core/n3494_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [25]),
	.I2(\top/processor/sha_core/w[59] [25]),
	.F(\top/processor/sha_core/n3494_178 )
);
defparam \top/processor/sha_core/n3494_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [24]),
	.I2(\top/processor/sha_core/w[3] [24]),
	.F(\top/processor/sha_core/n3495_172 )
);
defparam \top/processor/sha_core/n3495_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [24]),
	.I2(\top/processor/sha_core/w[11] [24]),
	.F(\top/processor/sha_core/n3495_173 )
);
defparam \top/processor/sha_core/n3495_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [24]),
	.I2(\top/processor/sha_core/w[19] [24]),
	.F(\top/processor/sha_core/n3495_174 )
);
defparam \top/processor/sha_core/n3495_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [24]),
	.I2(\top/processor/sha_core/w[27] [24]),
	.F(\top/processor/sha_core/n3495_175 )
);
defparam \top/processor/sha_core/n3495_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [31]),
	.I2(\top/processor/sha_core/w[43] [31]),
	.F(\top/processor/sha_core/n3488_172 )
);
defparam \top/processor/sha_core/n3488_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [24]),
	.I2(\top/processor/sha_core/w[35] [24]),
	.F(\top/processor/sha_core/n3495_176 )
);
defparam \top/processor/sha_core/n3495_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [24]),
	.I2(\top/processor/sha_core/w[43] [24]),
	.F(\top/processor/sha_core/n3495_177 )
);
defparam \top/processor/sha_core/n3495_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [24]),
	.I2(\top/processor/sha_core/w[51] [24]),
	.F(\top/processor/sha_core/n3495_178 )
);
defparam \top/processor/sha_core/n3495_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3495_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [24]),
	.I2(\top/processor/sha_core/w[59] [24]),
	.F(\top/processor/sha_core/n3495_179 )
);
defparam \top/processor/sha_core/n3495_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [23]),
	.I2(\top/processor/sha_core/w[3] [23]),
	.F(\top/processor/sha_core/n3496_172 )
);
defparam \top/processor/sha_core/n3496_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [23]),
	.I2(\top/processor/sha_core/w[11] [23]),
	.F(\top/processor/sha_core/n3496_173 )
);
defparam \top/processor/sha_core/n3496_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [23]),
	.I2(\top/processor/sha_core/w[19] [23]),
	.F(\top/processor/sha_core/n3496_174 )
);
defparam \top/processor/sha_core/n3496_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [23]),
	.I2(\top/processor/sha_core/w[27] [23]),
	.F(\top/processor/sha_core/n3496_175 )
);
defparam \top/processor/sha_core/n3496_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [23]),
	.I2(\top/processor/sha_core/w[35] [23]),
	.F(\top/processor/sha_core/n3496_176 )
);
defparam \top/processor/sha_core/n3496_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [23]),
	.I2(\top/processor/sha_core/w[43] [23]),
	.F(\top/processor/sha_core/n3496_177 )
);
defparam \top/processor/sha_core/n3496_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [31]),
	.I2(\top/processor/sha_core/w[51] [31]),
	.F(\top/processor/sha_core/n3488_173 )
);
defparam \top/processor/sha_core/n3488_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [23]),
	.I2(\top/processor/sha_core/w[51] [23]),
	.F(\top/processor/sha_core/n3496_178 )
);
defparam \top/processor/sha_core/n3496_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3496_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [23]),
	.I2(\top/processor/sha_core/w[59] [23]),
	.F(\top/processor/sha_core/n3496_179 )
);
defparam \top/processor/sha_core/n3496_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [22]),
	.I2(\top/processor/sha_core/w[3] [22]),
	.F(\top/processor/sha_core/n3497_172 )
);
defparam \top/processor/sha_core/n3497_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [22]),
	.I2(\top/processor/sha_core/w[11] [22]),
	.F(\top/processor/sha_core/n3497_173 )
);
defparam \top/processor/sha_core/n3497_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [22]),
	.I2(\top/processor/sha_core/w[19] [22]),
	.F(\top/processor/sha_core/n3497_174 )
);
defparam \top/processor/sha_core/n3497_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [22]),
	.I2(\top/processor/sha_core/w[27] [22]),
	.F(\top/processor/sha_core/n3497_175 )
);
defparam \top/processor/sha_core/n3497_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [22]),
	.I2(\top/processor/sha_core/w[35] [22]),
	.F(\top/processor/sha_core/n3497_176 )
);
defparam \top/processor/sha_core/n3497_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [22]),
	.I2(\top/processor/sha_core/w[43] [22]),
	.F(\top/processor/sha_core/n3497_177 )
);
defparam \top/processor/sha_core/n3497_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [22]),
	.I2(\top/processor/sha_core/w[51] [22]),
	.F(\top/processor/sha_core/n3497_178 )
);
defparam \top/processor/sha_core/n3497_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3497_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [22]),
	.I2(\top/processor/sha_core/w[59] [22]),
	.F(\top/processor/sha_core/n3497_179 )
);
defparam \top/processor/sha_core/n3497_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [31]),
	.I2(\top/processor/sha_core/w[59] [31]),
	.F(\top/processor/sha_core/n3488_174 )
);
defparam \top/processor/sha_core/n3488_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [21]),
	.I2(\top/processor/sha_core/w[3] [21]),
	.F(\top/processor/sha_core/n3498_172 )
);
defparam \top/processor/sha_core/n3498_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [21]),
	.I2(\top/processor/sha_core/w[11] [21]),
	.F(\top/processor/sha_core/n3498_173 )
);
defparam \top/processor/sha_core/n3498_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [21]),
	.I2(\top/processor/sha_core/w[19] [21]),
	.F(\top/processor/sha_core/n3498_174 )
);
defparam \top/processor/sha_core/n3498_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [21]),
	.I2(\top/processor/sha_core/w[27] [21]),
	.F(\top/processor/sha_core/n3498_175 )
);
defparam \top/processor/sha_core/n3498_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [21]),
	.I2(\top/processor/sha_core/w[35] [21]),
	.F(\top/processor/sha_core/n3498_176 )
);
defparam \top/processor/sha_core/n3498_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [21]),
	.I2(\top/processor/sha_core/w[43] [21]),
	.F(\top/processor/sha_core/n3498_177 )
);
defparam \top/processor/sha_core/n3498_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [21]),
	.I2(\top/processor/sha_core/w[51] [21]),
	.F(\top/processor/sha_core/n3498_178 )
);
defparam \top/processor/sha_core/n3498_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3498_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [21]),
	.I2(\top/processor/sha_core/w[59] [21]),
	.F(\top/processor/sha_core/n3498_179 )
);
defparam \top/processor/sha_core/n3498_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [20]),
	.I2(\top/processor/sha_core/w[3] [20]),
	.F(\top/processor/sha_core/n3499_172 )
);
defparam \top/processor/sha_core/n3499_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [20]),
	.I2(\top/processor/sha_core/w[11] [20]),
	.F(\top/processor/sha_core/n3499_173 )
);
defparam \top/processor/sha_core/n3499_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [30]),
	.I2(\top/processor/sha_core/w[3] [30]),
	.F(\top/processor/sha_core/n3489_172 )
);
defparam \top/processor/sha_core/n3489_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [20]),
	.I2(\top/processor/sha_core/w[19] [20]),
	.F(\top/processor/sha_core/n3499_174 )
);
defparam \top/processor/sha_core/n3499_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [20]),
	.I2(\top/processor/sha_core/w[27] [20]),
	.F(\top/processor/sha_core/n3499_175 )
);
defparam \top/processor/sha_core/n3499_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [20]),
	.I2(\top/processor/sha_core/w[35] [20]),
	.F(\top/processor/sha_core/n3499_176 )
);
defparam \top/processor/sha_core/n3499_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [20]),
	.I2(\top/processor/sha_core/w[43] [20]),
	.F(\top/processor/sha_core/n3499_177 )
);
defparam \top/processor/sha_core/n3499_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [20]),
	.I2(\top/processor/sha_core/w[51] [20]),
	.F(\top/processor/sha_core/n3499_178 )
);
defparam \top/processor/sha_core/n3499_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3499_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [20]),
	.I2(\top/processor/sha_core/w[59] [20]),
	.F(\top/processor/sha_core/n3499_179 )
);
defparam \top/processor/sha_core/n3499_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [19]),
	.I2(\top/processor/sha_core/w[3] [19]),
	.F(\top/processor/sha_core/n3500_172 )
);
defparam \top/processor/sha_core/n3500_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [19]),
	.I2(\top/processor/sha_core/w[11] [19]),
	.F(\top/processor/sha_core/n3500_173 )
);
defparam \top/processor/sha_core/n3500_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [19]),
	.I2(\top/processor/sha_core/w[19] [19]),
	.F(\top/processor/sha_core/n3500_174 )
);
defparam \top/processor/sha_core/n3500_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [19]),
	.I2(\top/processor/sha_core/w[27] [19]),
	.F(\top/processor/sha_core/n3500_175 )
);
defparam \top/processor/sha_core/n3500_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [30]),
	.I2(\top/processor/sha_core/w[11] [30]),
	.F(\top/processor/sha_core/n3489_173 )
);
defparam \top/processor/sha_core/n3489_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [31]),
	.I2(\top/processor/sha_core/w[3] [31]),
	.F(\top/processor/sha_core/n3488_175 )
);
defparam \top/processor/sha_core/n3488_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [19]),
	.I2(\top/processor/sha_core/w[35] [19]),
	.F(\top/processor/sha_core/n3500_176 )
);
defparam \top/processor/sha_core/n3500_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [19]),
	.I2(\top/processor/sha_core/w[43] [19]),
	.F(\top/processor/sha_core/n3500_177 )
);
defparam \top/processor/sha_core/n3500_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [19]),
	.I2(\top/processor/sha_core/w[51] [19]),
	.F(\top/processor/sha_core/n3500_178 )
);
defparam \top/processor/sha_core/n3500_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3500_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [19]),
	.I2(\top/processor/sha_core/w[59] [19]),
	.F(\top/processor/sha_core/n3500_179 )
);
defparam \top/processor/sha_core/n3500_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [18]),
	.I2(\top/processor/sha_core/w[3] [18]),
	.F(\top/processor/sha_core/n3501_172 )
);
defparam \top/processor/sha_core/n3501_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [18]),
	.I2(\top/processor/sha_core/w[11] [18]),
	.F(\top/processor/sha_core/n3501_173 )
);
defparam \top/processor/sha_core/n3501_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [18]),
	.I2(\top/processor/sha_core/w[19] [18]),
	.F(\top/processor/sha_core/n3501_174 )
);
defparam \top/processor/sha_core/n3501_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [18]),
	.I2(\top/processor/sha_core/w[27] [18]),
	.F(\top/processor/sha_core/n3501_175 )
);
defparam \top/processor/sha_core/n3501_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [18]),
	.I2(\top/processor/sha_core/w[35] [18]),
	.F(\top/processor/sha_core/n3501_176 )
);
defparam \top/processor/sha_core/n3501_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [18]),
	.I2(\top/processor/sha_core/w[43] [18]),
	.F(\top/processor/sha_core/n3501_177 )
);
defparam \top/processor/sha_core/n3501_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [30]),
	.I2(\top/processor/sha_core/w[19] [30]),
	.F(\top/processor/sha_core/n3489_174 )
);
defparam \top/processor/sha_core/n3489_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [18]),
	.I2(\top/processor/sha_core/w[51] [18]),
	.F(\top/processor/sha_core/n3501_178 )
);
defparam \top/processor/sha_core/n3501_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3501_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [18]),
	.I2(\top/processor/sha_core/w[59] [18]),
	.F(\top/processor/sha_core/n3501_179 )
);
defparam \top/processor/sha_core/n3501_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [17]),
	.I2(\top/processor/sha_core/w[3] [17]),
	.F(\top/processor/sha_core/n3502_172 )
);
defparam \top/processor/sha_core/n3502_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [17]),
	.I2(\top/processor/sha_core/w[11] [17]),
	.F(\top/processor/sha_core/n3502_173 )
);
defparam \top/processor/sha_core/n3502_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [17]),
	.I2(\top/processor/sha_core/w[19] [17]),
	.F(\top/processor/sha_core/n3502_174 )
);
defparam \top/processor/sha_core/n3502_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [17]),
	.I2(\top/processor/sha_core/w[27] [17]),
	.F(\top/processor/sha_core/n3502_175 )
);
defparam \top/processor/sha_core/n3502_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [17]),
	.I2(\top/processor/sha_core/w[35] [17]),
	.F(\top/processor/sha_core/n3502_176 )
);
defparam \top/processor/sha_core/n3502_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [17]),
	.I2(\top/processor/sha_core/w[43] [17]),
	.F(\top/processor/sha_core/n3502_177 )
);
defparam \top/processor/sha_core/n3502_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [17]),
	.I2(\top/processor/sha_core/w[51] [17]),
	.F(\top/processor/sha_core/n3502_178 )
);
defparam \top/processor/sha_core/n3502_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3502_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [17]),
	.I2(\top/processor/sha_core/w[59] [17]),
	.F(\top/processor/sha_core/n3502_179 )
);
defparam \top/processor/sha_core/n3502_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [30]),
	.I2(\top/processor/sha_core/w[27] [30]),
	.F(\top/processor/sha_core/n3489_175 )
);
defparam \top/processor/sha_core/n3489_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [16]),
	.I2(\top/processor/sha_core/w[3] [16]),
	.F(\top/processor/sha_core/n3503_172 )
);
defparam \top/processor/sha_core/n3503_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [16]),
	.I2(\top/processor/sha_core/w[11] [16]),
	.F(\top/processor/sha_core/n3503_173 )
);
defparam \top/processor/sha_core/n3503_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [16]),
	.I2(\top/processor/sha_core/w[19] [16]),
	.F(\top/processor/sha_core/n3503_174 )
);
defparam \top/processor/sha_core/n3503_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [16]),
	.I2(\top/processor/sha_core/w[27] [16]),
	.F(\top/processor/sha_core/n3503_175 )
);
defparam \top/processor/sha_core/n3503_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [16]),
	.I2(\top/processor/sha_core/w[35] [16]),
	.F(\top/processor/sha_core/n3503_176 )
);
defparam \top/processor/sha_core/n3503_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [16]),
	.I2(\top/processor/sha_core/w[43] [16]),
	.F(\top/processor/sha_core/n3503_177 )
);
defparam \top/processor/sha_core/n3503_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [16]),
	.I2(\top/processor/sha_core/w[51] [16]),
	.F(\top/processor/sha_core/n3503_178 )
);
defparam \top/processor/sha_core/n3503_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3503_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [16]),
	.I2(\top/processor/sha_core/w[59] [16]),
	.F(\top/processor/sha_core/n3503_179 )
);
defparam \top/processor/sha_core/n3503_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [15]),
	.I2(\top/processor/sha_core/w[3] [15]),
	.F(\top/processor/sha_core/n3504_172 )
);
defparam \top/processor/sha_core/n3504_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [15]),
	.I2(\top/processor/sha_core/w[11] [15]),
	.F(\top/processor/sha_core/n3504_173 )
);
defparam \top/processor/sha_core/n3504_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [30]),
	.I2(\top/processor/sha_core/w[35] [30]),
	.F(\top/processor/sha_core/n3489_176 )
);
defparam \top/processor/sha_core/n3489_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [15]),
	.I2(\top/processor/sha_core/w[19] [15]),
	.F(\top/processor/sha_core/n3504_174 )
);
defparam \top/processor/sha_core/n3504_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [15]),
	.I2(\top/processor/sha_core/w[27] [15]),
	.F(\top/processor/sha_core/n3504_175 )
);
defparam \top/processor/sha_core/n3504_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [15]),
	.I2(\top/processor/sha_core/w[35] [15]),
	.F(\top/processor/sha_core/n3504_176 )
);
defparam \top/processor/sha_core/n3504_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [15]),
	.I2(\top/processor/sha_core/w[43] [15]),
	.F(\top/processor/sha_core/n3504_177 )
);
defparam \top/processor/sha_core/n3504_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [15]),
	.I2(\top/processor/sha_core/w[51] [15]),
	.F(\top/processor/sha_core/n3504_178 )
);
defparam \top/processor/sha_core/n3504_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3504_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [15]),
	.I2(\top/processor/sha_core/w[59] [15]),
	.F(\top/processor/sha_core/n3504_179 )
);
defparam \top/processor/sha_core/n3504_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [14]),
	.I2(\top/processor/sha_core/w[3] [14]),
	.F(\top/processor/sha_core/n3505_172 )
);
defparam \top/processor/sha_core/n3505_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [14]),
	.I2(\top/processor/sha_core/w[11] [14]),
	.F(\top/processor/sha_core/n3505_173 )
);
defparam \top/processor/sha_core/n3505_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [14]),
	.I2(\top/processor/sha_core/w[19] [14]),
	.F(\top/processor/sha_core/n3505_174 )
);
defparam \top/processor/sha_core/n3505_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [14]),
	.I2(\top/processor/sha_core/w[27] [14]),
	.F(\top/processor/sha_core/n3505_175 )
);
defparam \top/processor/sha_core/n3505_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [30]),
	.I2(\top/processor/sha_core/w[43] [30]),
	.F(\top/processor/sha_core/n3489_177 )
);
defparam \top/processor/sha_core/n3489_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [14]),
	.I2(\top/processor/sha_core/w[35] [14]),
	.F(\top/processor/sha_core/n3505_176 )
);
defparam \top/processor/sha_core/n3505_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [14]),
	.I2(\top/processor/sha_core/w[43] [14]),
	.F(\top/processor/sha_core/n3505_177 )
);
defparam \top/processor/sha_core/n3505_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [14]),
	.I2(\top/processor/sha_core/w[51] [14]),
	.F(\top/processor/sha_core/n3505_178 )
);
defparam \top/processor/sha_core/n3505_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3505_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [14]),
	.I2(\top/processor/sha_core/w[59] [14]),
	.F(\top/processor/sha_core/n3505_179 )
);
defparam \top/processor/sha_core/n3505_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [13]),
	.I2(\top/processor/sha_core/w[3] [13]),
	.F(\top/processor/sha_core/n3506_172 )
);
defparam \top/processor/sha_core/n3506_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [13]),
	.I2(\top/processor/sha_core/w[11] [13]),
	.F(\top/processor/sha_core/n3506_173 )
);
defparam \top/processor/sha_core/n3506_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [13]),
	.I2(\top/processor/sha_core/w[19] [13]),
	.F(\top/processor/sha_core/n3506_174 )
);
defparam \top/processor/sha_core/n3506_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [13]),
	.I2(\top/processor/sha_core/w[27] [13]),
	.F(\top/processor/sha_core/n3506_175 )
);
defparam \top/processor/sha_core/n3506_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [13]),
	.I2(\top/processor/sha_core/w[35] [13]),
	.F(\top/processor/sha_core/n3506_176 )
);
defparam \top/processor/sha_core/n3506_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [13]),
	.I2(\top/processor/sha_core/w[43] [13]),
	.F(\top/processor/sha_core/n3506_177 )
);
defparam \top/processor/sha_core/n3506_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [30]),
	.I2(\top/processor/sha_core/w[51] [30]),
	.F(\top/processor/sha_core/n3489_178 )
);
defparam \top/processor/sha_core/n3489_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [13]),
	.I2(\top/processor/sha_core/w[51] [13]),
	.F(\top/processor/sha_core/n3506_178 )
);
defparam \top/processor/sha_core/n3506_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3506_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [13]),
	.I2(\top/processor/sha_core/w[59] [13]),
	.F(\top/processor/sha_core/n3506_179 )
);
defparam \top/processor/sha_core/n3506_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [12]),
	.I2(\top/processor/sha_core/w[3] [12]),
	.F(\top/processor/sha_core/n3507_172 )
);
defparam \top/processor/sha_core/n3507_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [12]),
	.I2(\top/processor/sha_core/w[11] [12]),
	.F(\top/processor/sha_core/n3507_173 )
);
defparam \top/processor/sha_core/n3507_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [12]),
	.I2(\top/processor/sha_core/w[19] [12]),
	.F(\top/processor/sha_core/n3507_174 )
);
defparam \top/processor/sha_core/n3507_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [12]),
	.I2(\top/processor/sha_core/w[27] [12]),
	.F(\top/processor/sha_core/n3507_175 )
);
defparam \top/processor/sha_core/n3507_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [12]),
	.I2(\top/processor/sha_core/w[35] [12]),
	.F(\top/processor/sha_core/n3507_176 )
);
defparam \top/processor/sha_core/n3507_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [12]),
	.I2(\top/processor/sha_core/w[43] [12]),
	.F(\top/processor/sha_core/n3507_177 )
);
defparam \top/processor/sha_core/n3507_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [12]),
	.I2(\top/processor/sha_core/w[51] [12]),
	.F(\top/processor/sha_core/n3507_178 )
);
defparam \top/processor/sha_core/n3507_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3507_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [12]),
	.I2(\top/processor/sha_core/w[59] [12]),
	.F(\top/processor/sha_core/n3507_179 )
);
defparam \top/processor/sha_core/n3507_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3489_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [30]),
	.I2(\top/processor/sha_core/w[59] [30]),
	.F(\top/processor/sha_core/n3489_179 )
);
defparam \top/processor/sha_core/n3489_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [11]),
	.I2(\top/processor/sha_core/w[3] [11]),
	.F(\top/processor/sha_core/n3508_172 )
);
defparam \top/processor/sha_core/n3508_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [11]),
	.I2(\top/processor/sha_core/w[11] [11]),
	.F(\top/processor/sha_core/n3508_173 )
);
defparam \top/processor/sha_core/n3508_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [11]),
	.I2(\top/processor/sha_core/w[19] [11]),
	.F(\top/processor/sha_core/n3508_174 )
);
defparam \top/processor/sha_core/n3508_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [11]),
	.I2(\top/processor/sha_core/w[27] [11]),
	.F(\top/processor/sha_core/n3508_175 )
);
defparam \top/processor/sha_core/n3508_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [11]),
	.I2(\top/processor/sha_core/w[35] [11]),
	.F(\top/processor/sha_core/n3508_176 )
);
defparam \top/processor/sha_core/n3508_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [11]),
	.I2(\top/processor/sha_core/w[43] [11]),
	.F(\top/processor/sha_core/n3508_177 )
);
defparam \top/processor/sha_core/n3508_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [11]),
	.I2(\top/processor/sha_core/w[51] [11]),
	.F(\top/processor/sha_core/n3508_178 )
);
defparam \top/processor/sha_core/n3508_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3508_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [11]),
	.I2(\top/processor/sha_core/w[59] [11]),
	.F(\top/processor/sha_core/n3508_179 )
);
defparam \top/processor/sha_core/n3508_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [10]),
	.I2(\top/processor/sha_core/w[3] [10]),
	.F(\top/processor/sha_core/n3509_172 )
);
defparam \top/processor/sha_core/n3509_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [10]),
	.I2(\top/processor/sha_core/w[11] [10]),
	.F(\top/processor/sha_core/n3509_173 )
);
defparam \top/processor/sha_core/n3509_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [29]),
	.I2(\top/processor/sha_core/w[3] [29]),
	.F(\top/processor/sha_core/n3490_172 )
);
defparam \top/processor/sha_core/n3490_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [10]),
	.I2(\top/processor/sha_core/w[19] [10]),
	.F(\top/processor/sha_core/n3509_174 )
);
defparam \top/processor/sha_core/n3509_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [10]),
	.I2(\top/processor/sha_core/w[27] [10]),
	.F(\top/processor/sha_core/n3509_175 )
);
defparam \top/processor/sha_core/n3509_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [10]),
	.I2(\top/processor/sha_core/w[35] [10]),
	.F(\top/processor/sha_core/n3509_176 )
);
defparam \top/processor/sha_core/n3509_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [10]),
	.I2(\top/processor/sha_core/w[43] [10]),
	.F(\top/processor/sha_core/n3509_177 )
);
defparam \top/processor/sha_core/n3509_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [10]),
	.I2(\top/processor/sha_core/w[51] [10]),
	.F(\top/processor/sha_core/n3509_178 )
);
defparam \top/processor/sha_core/n3509_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3509_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [10]),
	.I2(\top/processor/sha_core/w[59] [10]),
	.F(\top/processor/sha_core/n3509_179 )
);
defparam \top/processor/sha_core/n3509_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [9]),
	.I2(\top/processor/sha_core/w[3] [9]),
	.F(\top/processor/sha_core/n3510_172 )
);
defparam \top/processor/sha_core/n3510_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [9]),
	.I2(\top/processor/sha_core/w[11] [9]),
	.F(\top/processor/sha_core/n3510_173 )
);
defparam \top/processor/sha_core/n3510_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [9]),
	.I2(\top/processor/sha_core/w[19] [9]),
	.F(\top/processor/sha_core/n3510_174 )
);
defparam \top/processor/sha_core/n3510_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [9]),
	.I2(\top/processor/sha_core/w[27] [9]),
	.F(\top/processor/sha_core/n3510_175 )
);
defparam \top/processor/sha_core/n3510_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [29]),
	.I2(\top/processor/sha_core/w[11] [29]),
	.F(\top/processor/sha_core/n3490_173 )
);
defparam \top/processor/sha_core/n3490_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [9]),
	.I2(\top/processor/sha_core/w[35] [9]),
	.F(\top/processor/sha_core/n3510_176 )
);
defparam \top/processor/sha_core/n3510_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [9]),
	.I2(\top/processor/sha_core/w[43] [9]),
	.F(\top/processor/sha_core/n3510_177 )
);
defparam \top/processor/sha_core/n3510_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [9]),
	.I2(\top/processor/sha_core/w[51] [9]),
	.F(\top/processor/sha_core/n3510_178 )
);
defparam \top/processor/sha_core/n3510_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3510_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [9]),
	.I2(\top/processor/sha_core/w[59] [9]),
	.F(\top/processor/sha_core/n3510_179 )
);
defparam \top/processor/sha_core/n3510_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [8]),
	.I2(\top/processor/sha_core/w[3] [8]),
	.F(\top/processor/sha_core/n3511_172 )
);
defparam \top/processor/sha_core/n3511_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [8]),
	.I2(\top/processor/sha_core/w[11] [8]),
	.F(\top/processor/sha_core/n3511_173 )
);
defparam \top/processor/sha_core/n3511_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [8]),
	.I2(\top/processor/sha_core/w[19] [8]),
	.F(\top/processor/sha_core/n3511_174 )
);
defparam \top/processor/sha_core/n3511_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [8]),
	.I2(\top/processor/sha_core/w[27] [8]),
	.F(\top/processor/sha_core/n3511_175 )
);
defparam \top/processor/sha_core/n3511_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [8]),
	.I2(\top/processor/sha_core/w[35] [8]),
	.F(\top/processor/sha_core/n3511_176 )
);
defparam \top/processor/sha_core/n3511_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [8]),
	.I2(\top/processor/sha_core/w[43] [8]),
	.F(\top/processor/sha_core/n3511_177 )
);
defparam \top/processor/sha_core/n3511_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [29]),
	.I2(\top/processor/sha_core/w[19] [29]),
	.F(\top/processor/sha_core/n3490_174 )
);
defparam \top/processor/sha_core/n3490_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [8]),
	.I2(\top/processor/sha_core/w[51] [8]),
	.F(\top/processor/sha_core/n3511_178 )
);
defparam \top/processor/sha_core/n3511_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3511_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [8]),
	.I2(\top/processor/sha_core/w[59] [8]),
	.F(\top/processor/sha_core/n3511_179 )
);
defparam \top/processor/sha_core/n3511_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [7]),
	.I2(\top/processor/sha_core/w[3] [7]),
	.F(\top/processor/sha_core/n3512_172 )
);
defparam \top/processor/sha_core/n3512_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [7]),
	.I2(\top/processor/sha_core/w[11] [7]),
	.F(\top/processor/sha_core/n3512_173 )
);
defparam \top/processor/sha_core/n3512_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [7]),
	.I2(\top/processor/sha_core/w[19] [7]),
	.F(\top/processor/sha_core/n3512_174 )
);
defparam \top/processor/sha_core/n3512_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [7]),
	.I2(\top/processor/sha_core/w[27] [7]),
	.F(\top/processor/sha_core/n3512_175 )
);
defparam \top/processor/sha_core/n3512_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [7]),
	.I2(\top/processor/sha_core/w[35] [7]),
	.F(\top/processor/sha_core/n3512_176 )
);
defparam \top/processor/sha_core/n3512_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [7]),
	.I2(\top/processor/sha_core/w[43] [7]),
	.F(\top/processor/sha_core/n3512_177 )
);
defparam \top/processor/sha_core/n3512_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [7]),
	.I2(\top/processor/sha_core/w[51] [7]),
	.F(\top/processor/sha_core/n3512_178 )
);
defparam \top/processor/sha_core/n3512_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3512_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [7]),
	.I2(\top/processor/sha_core/w[59] [7]),
	.F(\top/processor/sha_core/n3512_179 )
);
defparam \top/processor/sha_core/n3512_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [29]),
	.I2(\top/processor/sha_core/w[27] [29]),
	.F(\top/processor/sha_core/n3490_175 )
);
defparam \top/processor/sha_core/n3490_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [31]),
	.I2(\top/processor/sha_core/w[11] [31]),
	.F(\top/processor/sha_core/n3488_176 )
);
defparam \top/processor/sha_core/n3488_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [6]),
	.I2(\top/processor/sha_core/w[3] [6]),
	.F(\top/processor/sha_core/n3513_172 )
);
defparam \top/processor/sha_core/n3513_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [6]),
	.I2(\top/processor/sha_core/w[11] [6]),
	.F(\top/processor/sha_core/n3513_173 )
);
defparam \top/processor/sha_core/n3513_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [6]),
	.I2(\top/processor/sha_core/w[19] [6]),
	.F(\top/processor/sha_core/n3513_174 )
);
defparam \top/processor/sha_core/n3513_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [6]),
	.I2(\top/processor/sha_core/w[27] [6]),
	.F(\top/processor/sha_core/n3513_175 )
);
defparam \top/processor/sha_core/n3513_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [6]),
	.I2(\top/processor/sha_core/w[35] [6]),
	.F(\top/processor/sha_core/n3513_176 )
);
defparam \top/processor/sha_core/n3513_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [6]),
	.I2(\top/processor/sha_core/w[43] [6]),
	.F(\top/processor/sha_core/n3513_177 )
);
defparam \top/processor/sha_core/n3513_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [6]),
	.I2(\top/processor/sha_core/w[51] [6]),
	.F(\top/processor/sha_core/n3513_178 )
);
defparam \top/processor/sha_core/n3513_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3513_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [6]),
	.I2(\top/processor/sha_core/w[59] [6]),
	.F(\top/processor/sha_core/n3513_179 )
);
defparam \top/processor/sha_core/n3513_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [5]),
	.I2(\top/processor/sha_core/w[3] [5]),
	.F(\top/processor/sha_core/n3514_172 )
);
defparam \top/processor/sha_core/n3514_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [5]),
	.I2(\top/processor/sha_core/w[11] [5]),
	.F(\top/processor/sha_core/n3514_173 )
);
defparam \top/processor/sha_core/n3514_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [29]),
	.I2(\top/processor/sha_core/w[35] [29]),
	.F(\top/processor/sha_core/n3490_176 )
);
defparam \top/processor/sha_core/n3490_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [5]),
	.I2(\top/processor/sha_core/w[19] [5]),
	.F(\top/processor/sha_core/n3514_174 )
);
defparam \top/processor/sha_core/n3514_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [5]),
	.I2(\top/processor/sha_core/w[27] [5]),
	.F(\top/processor/sha_core/n3514_175 )
);
defparam \top/processor/sha_core/n3514_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [5]),
	.I2(\top/processor/sha_core/w[35] [5]),
	.F(\top/processor/sha_core/n3514_176 )
);
defparam \top/processor/sha_core/n3514_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [5]),
	.I2(\top/processor/sha_core/w[43] [5]),
	.F(\top/processor/sha_core/n3514_177 )
);
defparam \top/processor/sha_core/n3514_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [5]),
	.I2(\top/processor/sha_core/w[51] [5]),
	.F(\top/processor/sha_core/n3514_178 )
);
defparam \top/processor/sha_core/n3514_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3514_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [5]),
	.I2(\top/processor/sha_core/w[59] [5]),
	.F(\top/processor/sha_core/n3514_179 )
);
defparam \top/processor/sha_core/n3514_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [4]),
	.I2(\top/processor/sha_core/w[3] [4]),
	.F(\top/processor/sha_core/n3515_172 )
);
defparam \top/processor/sha_core/n3515_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [4]),
	.I2(\top/processor/sha_core/w[11] [4]),
	.F(\top/processor/sha_core/n3515_173 )
);
defparam \top/processor/sha_core/n3515_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [4]),
	.I2(\top/processor/sha_core/w[19] [4]),
	.F(\top/processor/sha_core/n3515_174 )
);
defparam \top/processor/sha_core/n3515_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [4]),
	.I2(\top/processor/sha_core/w[27] [4]),
	.F(\top/processor/sha_core/n3515_175 )
);
defparam \top/processor/sha_core/n3515_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [29]),
	.I2(\top/processor/sha_core/w[43] [29]),
	.F(\top/processor/sha_core/n3490_177 )
);
defparam \top/processor/sha_core/n3490_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [4]),
	.I2(\top/processor/sha_core/w[35] [4]),
	.F(\top/processor/sha_core/n3515_176 )
);
defparam \top/processor/sha_core/n3515_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [4]),
	.I2(\top/processor/sha_core/w[43] [4]),
	.F(\top/processor/sha_core/n3515_177 )
);
defparam \top/processor/sha_core/n3515_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [4]),
	.I2(\top/processor/sha_core/w[51] [4]),
	.F(\top/processor/sha_core/n3515_178 )
);
defparam \top/processor/sha_core/n3515_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3515_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [4]),
	.I2(\top/processor/sha_core/w[59] [4]),
	.F(\top/processor/sha_core/n3515_179 )
);
defparam \top/processor/sha_core/n3515_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [3]),
	.I2(\top/processor/sha_core/w[3] [3]),
	.F(\top/processor/sha_core/n3516_172 )
);
defparam \top/processor/sha_core/n3516_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [3]),
	.I2(\top/processor/sha_core/w[11] [3]),
	.F(\top/processor/sha_core/n3516_173 )
);
defparam \top/processor/sha_core/n3516_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [3]),
	.I2(\top/processor/sha_core/w[19] [3]),
	.F(\top/processor/sha_core/n3516_174 )
);
defparam \top/processor/sha_core/n3516_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [3]),
	.I2(\top/processor/sha_core/w[27] [3]),
	.F(\top/processor/sha_core/n3516_175 )
);
defparam \top/processor/sha_core/n3516_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [3]),
	.I2(\top/processor/sha_core/w[35] [3]),
	.F(\top/processor/sha_core/n3516_176 )
);
defparam \top/processor/sha_core/n3516_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [3]),
	.I2(\top/processor/sha_core/w[43] [3]),
	.F(\top/processor/sha_core/n3516_177 )
);
defparam \top/processor/sha_core/n3516_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [29]),
	.I2(\top/processor/sha_core/w[51] [29]),
	.F(\top/processor/sha_core/n3490_178 )
);
defparam \top/processor/sha_core/n3490_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [3]),
	.I2(\top/processor/sha_core/w[51] [3]),
	.F(\top/processor/sha_core/n3516_178 )
);
defparam \top/processor/sha_core/n3516_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3516_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [3]),
	.I2(\top/processor/sha_core/w[59] [3]),
	.F(\top/processor/sha_core/n3516_179 )
);
defparam \top/processor/sha_core/n3516_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [2]),
	.I2(\top/processor/sha_core/w[3] [2]),
	.F(\top/processor/sha_core/n3517_172 )
);
defparam \top/processor/sha_core/n3517_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [2]),
	.I2(\top/processor/sha_core/w[11] [2]),
	.F(\top/processor/sha_core/n3517_173 )
);
defparam \top/processor/sha_core/n3517_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [2]),
	.I2(\top/processor/sha_core/w[19] [2]),
	.F(\top/processor/sha_core/n3517_174 )
);
defparam \top/processor/sha_core/n3517_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [2]),
	.I2(\top/processor/sha_core/w[27] [2]),
	.F(\top/processor/sha_core/n3517_175 )
);
defparam \top/processor/sha_core/n3517_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [2]),
	.I2(\top/processor/sha_core/w[35] [2]),
	.F(\top/processor/sha_core/n3517_176 )
);
defparam \top/processor/sha_core/n3517_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [2]),
	.I2(\top/processor/sha_core/w[43] [2]),
	.F(\top/processor/sha_core/n3517_177 )
);
defparam \top/processor/sha_core/n3517_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [2]),
	.I2(\top/processor/sha_core/w[51] [2]),
	.F(\top/processor/sha_core/n3517_178 )
);
defparam \top/processor/sha_core/n3517_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3517_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [2]),
	.I2(\top/processor/sha_core/w[59] [2]),
	.F(\top/processor/sha_core/n3517_179 )
);
defparam \top/processor/sha_core/n3517_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3490_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [29]),
	.I2(\top/processor/sha_core/w[59] [29]),
	.F(\top/processor/sha_core/n3490_179 )
);
defparam \top/processor/sha_core/n3490_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [1]),
	.I2(\top/processor/sha_core/w[3] [1]),
	.F(\top/processor/sha_core/n3518_172 )
);
defparam \top/processor/sha_core/n3518_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [1]),
	.I2(\top/processor/sha_core/w[11] [1]),
	.F(\top/processor/sha_core/n3518_173 )
);
defparam \top/processor/sha_core/n3518_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [1]),
	.I2(\top/processor/sha_core/w[19] [1]),
	.F(\top/processor/sha_core/n3518_174 )
);
defparam \top/processor/sha_core/n3518_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [1]),
	.I2(\top/processor/sha_core/w[27] [1]),
	.F(\top/processor/sha_core/n3518_175 )
);
defparam \top/processor/sha_core/n3518_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [1]),
	.I2(\top/processor/sha_core/w[35] [1]),
	.F(\top/processor/sha_core/n3518_176 )
);
defparam \top/processor/sha_core/n3518_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [1]),
	.I2(\top/processor/sha_core/w[43] [1]),
	.F(\top/processor/sha_core/n3518_177 )
);
defparam \top/processor/sha_core/n3518_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [1]),
	.I2(\top/processor/sha_core/w[51] [1]),
	.F(\top/processor/sha_core/n3518_178 )
);
defparam \top/processor/sha_core/n3518_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3518_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [1]),
	.I2(\top/processor/sha_core/w[59] [1]),
	.F(\top/processor/sha_core/n3518_179 )
);
defparam \top/processor/sha_core/n3518_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [0]),
	.I2(\top/processor/sha_core/w[3] [0]),
	.F(\top/processor/sha_core/n3519_172 )
);
defparam \top/processor/sha_core/n3519_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [0]),
	.I2(\top/processor/sha_core/w[11] [0]),
	.F(\top/processor/sha_core/n3519_173 )
);
defparam \top/processor/sha_core/n3519_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [28]),
	.I2(\top/processor/sha_core/w[3] [28]),
	.F(\top/processor/sha_core/n3491_172 )
);
defparam \top/processor/sha_core/n3491_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [0]),
	.I2(\top/processor/sha_core/w[19] [0]),
	.F(\top/processor/sha_core/n3519_174 )
);
defparam \top/processor/sha_core/n3519_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [0]),
	.I2(\top/processor/sha_core/w[27] [0]),
	.F(\top/processor/sha_core/n3519_175 )
);
defparam \top/processor/sha_core/n3519_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [0]),
	.I2(\top/processor/sha_core/w[35] [0]),
	.F(\top/processor/sha_core/n3519_176 )
);
defparam \top/processor/sha_core/n3519_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [0]),
	.I2(\top/processor/sha_core/w[43] [0]),
	.F(\top/processor/sha_core/n3519_177 )
);
defparam \top/processor/sha_core/n3519_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [0]),
	.I2(\top/processor/sha_core/w[51] [0]),
	.F(\top/processor/sha_core/n3519_178 )
);
defparam \top/processor/sha_core/n3519_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3519_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [0]),
	.I2(\top/processor/sha_core/w[59] [0]),
	.F(\top/processor/sha_core/n3519_179 )
);
defparam \top/processor/sha_core/n3519_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [28]),
	.I2(\top/processor/sha_core/w[11] [28]),
	.F(\top/processor/sha_core/n3491_173 )
);
defparam \top/processor/sha_core/n3491_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [28]),
	.I2(\top/processor/sha_core/w[19] [28]),
	.F(\top/processor/sha_core/n3491_174 )
);
defparam \top/processor/sha_core/n3491_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [28]),
	.I2(\top/processor/sha_core/w[27] [28]),
	.F(\top/processor/sha_core/n3491_175 )
);
defparam \top/processor/sha_core/n3491_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [28]),
	.I2(\top/processor/sha_core/w[35] [28]),
	.F(\top/processor/sha_core/n3491_176 )
);
defparam \top/processor/sha_core/n3491_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [28]),
	.I2(\top/processor/sha_core/w[43] [28]),
	.F(\top/processor/sha_core/n3491_177 )
);
defparam \top/processor/sha_core/n3491_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [31]),
	.I2(\top/processor/sha_core/w[19] [31]),
	.F(\top/processor/sha_core/n3488_177 )
);
defparam \top/processor/sha_core/n3488_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [28]),
	.I2(\top/processor/sha_core/w[51] [28]),
	.F(\top/processor/sha_core/n3491_178 )
);
defparam \top/processor/sha_core/n3491_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3491_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [28]),
	.I2(\top/processor/sha_core/w[59] [28]),
	.F(\top/processor/sha_core/n3491_179 )
);
defparam \top/processor/sha_core/n3491_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [27]),
	.I2(\top/processor/sha_core/w[3] [27]),
	.F(\top/processor/sha_core/n3492_172 )
);
defparam \top/processor/sha_core/n3492_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [27]),
	.I2(\top/processor/sha_core/w[11] [27]),
	.F(\top/processor/sha_core/n3492_173 )
);
defparam \top/processor/sha_core/n3492_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [27]),
	.I2(\top/processor/sha_core/w[19] [27]),
	.F(\top/processor/sha_core/n3492_174 )
);
defparam \top/processor/sha_core/n3492_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [27]),
	.I2(\top/processor/sha_core/w[27] [27]),
	.F(\top/processor/sha_core/n3492_175 )
);
defparam \top/processor/sha_core/n3492_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [27]),
	.I2(\top/processor/sha_core/w[35] [27]),
	.F(\top/processor/sha_core/n3492_176 )
);
defparam \top/processor/sha_core/n3492_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [27]),
	.I2(\top/processor/sha_core/w[43] [27]),
	.F(\top/processor/sha_core/n3492_177 )
);
defparam \top/processor/sha_core/n3492_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [27]),
	.I2(\top/processor/sha_core/w[51] [27]),
	.F(\top/processor/sha_core/n3492_178 )
);
defparam \top/processor/sha_core/n3492_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3492_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [27]),
	.I2(\top/processor/sha_core/w[59] [27]),
	.F(\top/processor/sha_core/n3492_179 )
);
defparam \top/processor/sha_core/n3492_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [31]),
	.I2(\top/processor/sha_core/w[27] [31]),
	.F(\top/processor/sha_core/n3488_178 )
);
defparam \top/processor/sha_core/n3488_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s159  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [26]),
	.I2(\top/processor/sha_core/w[3] [26]),
	.F(\top/processor/sha_core/n3493_172 )
);
defparam \top/processor/sha_core/n3493_s159 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s160  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [26]),
	.I2(\top/processor/sha_core/w[11] [26]),
	.F(\top/processor/sha_core/n3493_173 )
);
defparam \top/processor/sha_core/n3493_s160 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s161  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[18] [26]),
	.I2(\top/processor/sha_core/w[19] [26]),
	.F(\top/processor/sha_core/n3493_174 )
);
defparam \top/processor/sha_core/n3493_s161 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s162  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[26] [26]),
	.I2(\top/processor/sha_core/w[27] [26]),
	.F(\top/processor/sha_core/n3493_175 )
);
defparam \top/processor/sha_core/n3493_s162 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s163  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[34] [26]),
	.I2(\top/processor/sha_core/w[35] [26]),
	.F(\top/processor/sha_core/n3493_176 )
);
defparam \top/processor/sha_core/n3493_s163 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s164  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[42] [26]),
	.I2(\top/processor/sha_core/w[43] [26]),
	.F(\top/processor/sha_core/n3493_177 )
);
defparam \top/processor/sha_core/n3493_s164 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[50] [26]),
	.I2(\top/processor/sha_core/w[51] [26]),
	.F(\top/processor/sha_core/n3493_178 )
);
defparam \top/processor/sha_core/n3493_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3493_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[58] [26]),
	.I2(\top/processor/sha_core/w[59] [26]),
	.F(\top/processor/sha_core/n3493_179 )
);
defparam \top/processor/sha_core/n3493_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s165  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[2] [25]),
	.I2(\top/processor/sha_core/w[3] [25]),
	.F(\top/processor/sha_core/n3494_179 )
);
defparam \top/processor/sha_core/n3494_s165 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3494_s166  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/w[10] [25]),
	.I2(\top/processor/sha_core/w[11] [25]),
	.F(\top/processor/sha_core/n3494_180 )
);
defparam \top/processor/sha_core/n3494_s166 .INIT=8'hE4;
LUT3 \top/processor/sha_core/n3488_s166  (
	.I0(\top/processor/sha_core/w[34] [31]),
	.I1(\top/processor/sha_core/w[35] [31]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.F(\top/processor/sha_core/n3488_179 )
);
defparam \top/processor/sha_core/n3488_s166 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s218  (
	.I0(\top/processor/sha_core/w[0] [31]),
	.I1(\top/processor/sha_core/w[1] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_132 )
);
defparam \top/processor/sha_core/n327_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s219  (
	.I0(\top/processor/sha_core/w[2] [31]),
	.I1(\top/processor/sha_core/w[3] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_133 )
);
defparam \top/processor/sha_core/n327_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s220  (
	.I0(\top/processor/sha_core/w[4] [31]),
	.I1(\top/processor/sha_core/w[5] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_134 )
);
defparam \top/processor/sha_core/n327_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s221  (
	.I0(\top/processor/sha_core/w[6] [31]),
	.I1(\top/processor/sha_core/w[7] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_135 )
);
defparam \top/processor/sha_core/n327_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s222  (
	.I0(\top/processor/sha_core/w[8] [31]),
	.I1(\top/processor/sha_core/w[9] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_136 )
);
defparam \top/processor/sha_core/n327_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s223  (
	.I0(\top/processor/sha_core/w[10] [31]),
	.I1(\top/processor/sha_core/w[11] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_137 )
);
defparam \top/processor/sha_core/n327_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s224  (
	.I0(\top/processor/sha_core/w[12] [31]),
	.I1(\top/processor/sha_core/w[13] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_138 )
);
defparam \top/processor/sha_core/n327_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s225  (
	.I0(\top/processor/sha_core/w[14] [31]),
	.I1(\top/processor/sha_core/w[15] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_139 )
);
defparam \top/processor/sha_core/n327_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s226  (
	.I0(\top/processor/sha_core/w[16] [31]),
	.I1(\top/processor/sha_core/w[17] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_140 )
);
defparam \top/processor/sha_core/n327_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s227  (
	.I0(\top/processor/sha_core/w[18] [31]),
	.I1(\top/processor/sha_core/w[19] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_141 )
);
defparam \top/processor/sha_core/n327_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s228  (
	.I0(\top/processor/sha_core/w[20] [31]),
	.I1(\top/processor/sha_core/w[21] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_142 )
);
defparam \top/processor/sha_core/n327_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s229  (
	.I0(\top/processor/sha_core/w[22] [31]),
	.I1(\top/processor/sha_core/w[23] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_143 )
);
defparam \top/processor/sha_core/n327_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s230  (
	.I0(\top/processor/sha_core/w[24] [31]),
	.I1(\top/processor/sha_core/w[25] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_144 )
);
defparam \top/processor/sha_core/n327_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s231  (
	.I0(\top/processor/sha_core/w[26] [31]),
	.I1(\top/processor/sha_core/w[27] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_145 )
);
defparam \top/processor/sha_core/n327_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s232  (
	.I0(\top/processor/sha_core/w[28] [31]),
	.I1(\top/processor/sha_core/w[29] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_146 )
);
defparam \top/processor/sha_core/n327_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s233  (
	.I0(\top/processor/sha_core/w[30] [31]),
	.I1(\top/processor/sha_core/w[31] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_147 )
);
defparam \top/processor/sha_core/n327_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s234  (
	.I0(\top/processor/sha_core/w[32] [31]),
	.I1(\top/processor/sha_core/w[33] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_148 )
);
defparam \top/processor/sha_core/n327_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s235  (
	.I0(\top/processor/sha_core/w[34] [31]),
	.I1(\top/processor/sha_core/w[35] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_149 )
);
defparam \top/processor/sha_core/n327_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s236  (
	.I0(\top/processor/sha_core/w[36] [31]),
	.I1(\top/processor/sha_core/w[37] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_150 )
);
defparam \top/processor/sha_core/n327_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s237  (
	.I0(\top/processor/sha_core/w[38] [31]),
	.I1(\top/processor/sha_core/w[39] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_151 )
);
defparam \top/processor/sha_core/n327_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s238  (
	.I0(\top/processor/sha_core/w[40] [31]),
	.I1(\top/processor/sha_core/w[41] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_152 )
);
defparam \top/processor/sha_core/n327_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s239  (
	.I0(\top/processor/sha_core/w[42] [31]),
	.I1(\top/processor/sha_core/w[43] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_153 )
);
defparam \top/processor/sha_core/n327_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s240  (
	.I0(\top/processor/sha_core/w[44] [31]),
	.I1(\top/processor/sha_core/w[45] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_154 )
);
defparam \top/processor/sha_core/n327_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s241  (
	.I0(\top/processor/sha_core/w[46] [31]),
	.I1(\top/processor/sha_core/w[47] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_155 )
);
defparam \top/processor/sha_core/n327_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s242  (
	.I0(\top/processor/sha_core/w[48] [31]),
	.I1(\top/processor/sha_core/w[49] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_156 )
);
defparam \top/processor/sha_core/n327_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s243  (
	.I0(\top/processor/sha_core/w[50] [31]),
	.I1(\top/processor/sha_core/w[51] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_157 )
);
defparam \top/processor/sha_core/n327_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s244  (
	.I0(\top/processor/sha_core/w[52] [31]),
	.I1(\top/processor/sha_core/w[53] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_158 )
);
defparam \top/processor/sha_core/n327_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s245  (
	.I0(\top/processor/sha_core/w[54] [31]),
	.I1(\top/processor/sha_core/w[55] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_159 )
);
defparam \top/processor/sha_core/n327_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s246  (
	.I0(\top/processor/sha_core/w[56] [31]),
	.I1(\top/processor/sha_core/w[57] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_160 )
);
defparam \top/processor/sha_core/n327_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s247  (
	.I0(\top/processor/sha_core/w[58] [31]),
	.I1(\top/processor/sha_core/w[59] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_161 )
);
defparam \top/processor/sha_core/n327_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s248  (
	.I0(\top/processor/sha_core/w[60] [31]),
	.I1(\top/processor/sha_core/w[61] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_162 )
);
defparam \top/processor/sha_core/n327_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n327_s249  (
	.I0(\top/processor/sha_core/w[62] [31]),
	.I1(\top/processor/sha_core/w[63] [31]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n327_163 )
);
defparam \top/processor/sha_core/n327_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s218  (
	.I0(\top/processor/sha_core/w[0] [30]),
	.I1(\top/processor/sha_core/w[1] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_132 )
);
defparam \top/processor/sha_core/n328_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s219  (
	.I0(\top/processor/sha_core/w[2] [30]),
	.I1(\top/processor/sha_core/w[3] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_133 )
);
defparam \top/processor/sha_core/n328_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s220  (
	.I0(\top/processor/sha_core/w[4] [30]),
	.I1(\top/processor/sha_core/w[5] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_134 )
);
defparam \top/processor/sha_core/n328_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s221  (
	.I0(\top/processor/sha_core/w[6] [30]),
	.I1(\top/processor/sha_core/w[7] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_135 )
);
defparam \top/processor/sha_core/n328_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s222  (
	.I0(\top/processor/sha_core/w[8] [30]),
	.I1(\top/processor/sha_core/w[9] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_136 )
);
defparam \top/processor/sha_core/n328_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s223  (
	.I0(\top/processor/sha_core/w[10] [30]),
	.I1(\top/processor/sha_core/w[11] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_137 )
);
defparam \top/processor/sha_core/n328_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s224  (
	.I0(\top/processor/sha_core/w[12] [30]),
	.I1(\top/processor/sha_core/w[13] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_138 )
);
defparam \top/processor/sha_core/n328_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s225  (
	.I0(\top/processor/sha_core/w[14] [30]),
	.I1(\top/processor/sha_core/w[15] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_139 )
);
defparam \top/processor/sha_core/n328_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s226  (
	.I0(\top/processor/sha_core/w[16] [30]),
	.I1(\top/processor/sha_core/w[17] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_140 )
);
defparam \top/processor/sha_core/n328_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s227  (
	.I0(\top/processor/sha_core/w[18] [30]),
	.I1(\top/processor/sha_core/w[19] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_141 )
);
defparam \top/processor/sha_core/n328_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s228  (
	.I0(\top/processor/sha_core/w[20] [30]),
	.I1(\top/processor/sha_core/w[21] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_142 )
);
defparam \top/processor/sha_core/n328_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s229  (
	.I0(\top/processor/sha_core/w[22] [30]),
	.I1(\top/processor/sha_core/w[23] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_143 )
);
defparam \top/processor/sha_core/n328_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s230  (
	.I0(\top/processor/sha_core/w[24] [30]),
	.I1(\top/processor/sha_core/w[25] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_144 )
);
defparam \top/processor/sha_core/n328_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s231  (
	.I0(\top/processor/sha_core/w[26] [30]),
	.I1(\top/processor/sha_core/w[27] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_145 )
);
defparam \top/processor/sha_core/n328_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s232  (
	.I0(\top/processor/sha_core/w[28] [30]),
	.I1(\top/processor/sha_core/w[29] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_146 )
);
defparam \top/processor/sha_core/n328_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s233  (
	.I0(\top/processor/sha_core/w[30] [30]),
	.I1(\top/processor/sha_core/w[31] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_147 )
);
defparam \top/processor/sha_core/n328_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s234  (
	.I0(\top/processor/sha_core/w[32] [30]),
	.I1(\top/processor/sha_core/w[33] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_148 )
);
defparam \top/processor/sha_core/n328_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s235  (
	.I0(\top/processor/sha_core/w[34] [30]),
	.I1(\top/processor/sha_core/w[35] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_149 )
);
defparam \top/processor/sha_core/n328_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s236  (
	.I0(\top/processor/sha_core/w[36] [30]),
	.I1(\top/processor/sha_core/w[37] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_150 )
);
defparam \top/processor/sha_core/n328_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s237  (
	.I0(\top/processor/sha_core/w[38] [30]),
	.I1(\top/processor/sha_core/w[39] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_151 )
);
defparam \top/processor/sha_core/n328_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s238  (
	.I0(\top/processor/sha_core/w[40] [30]),
	.I1(\top/processor/sha_core/w[41] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_152 )
);
defparam \top/processor/sha_core/n328_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s239  (
	.I0(\top/processor/sha_core/w[42] [30]),
	.I1(\top/processor/sha_core/w[43] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_153 )
);
defparam \top/processor/sha_core/n328_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s240  (
	.I0(\top/processor/sha_core/w[44] [30]),
	.I1(\top/processor/sha_core/w[45] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_154 )
);
defparam \top/processor/sha_core/n328_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s241  (
	.I0(\top/processor/sha_core/w[46] [30]),
	.I1(\top/processor/sha_core/w[47] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_155 )
);
defparam \top/processor/sha_core/n328_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s242  (
	.I0(\top/processor/sha_core/w[48] [30]),
	.I1(\top/processor/sha_core/w[49] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_156 )
);
defparam \top/processor/sha_core/n328_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s243  (
	.I0(\top/processor/sha_core/w[50] [30]),
	.I1(\top/processor/sha_core/w[51] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_157 )
);
defparam \top/processor/sha_core/n328_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s244  (
	.I0(\top/processor/sha_core/w[52] [30]),
	.I1(\top/processor/sha_core/w[53] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_158 )
);
defparam \top/processor/sha_core/n328_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s245  (
	.I0(\top/processor/sha_core/w[54] [30]),
	.I1(\top/processor/sha_core/w[55] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_159 )
);
defparam \top/processor/sha_core/n328_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s246  (
	.I0(\top/processor/sha_core/w[56] [30]),
	.I1(\top/processor/sha_core/w[57] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_160 )
);
defparam \top/processor/sha_core/n328_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s247  (
	.I0(\top/processor/sha_core/w[58] [30]),
	.I1(\top/processor/sha_core/w[59] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_161 )
);
defparam \top/processor/sha_core/n328_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s248  (
	.I0(\top/processor/sha_core/w[60] [30]),
	.I1(\top/processor/sha_core/w[61] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_162 )
);
defparam \top/processor/sha_core/n328_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s249  (
	.I0(\top/processor/sha_core/w[62] [30]),
	.I1(\top/processor/sha_core/w[63] [30]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n328_163 )
);
defparam \top/processor/sha_core/n328_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s218  (
	.I0(\top/processor/sha_core/w[0] [29]),
	.I1(\top/processor/sha_core/w[1] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_132 )
);
defparam \top/processor/sha_core/n329_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s219  (
	.I0(\top/processor/sha_core/w[2] [29]),
	.I1(\top/processor/sha_core/w[3] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_133 )
);
defparam \top/processor/sha_core/n329_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s220  (
	.I0(\top/processor/sha_core/w[4] [29]),
	.I1(\top/processor/sha_core/w[5] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_134 )
);
defparam \top/processor/sha_core/n329_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s221  (
	.I0(\top/processor/sha_core/w[6] [29]),
	.I1(\top/processor/sha_core/w[7] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_135 )
);
defparam \top/processor/sha_core/n329_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s222  (
	.I0(\top/processor/sha_core/w[8] [29]),
	.I1(\top/processor/sha_core/w[9] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_136 )
);
defparam \top/processor/sha_core/n329_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s223  (
	.I0(\top/processor/sha_core/w[10] [29]),
	.I1(\top/processor/sha_core/w[11] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_137 )
);
defparam \top/processor/sha_core/n329_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s224  (
	.I0(\top/processor/sha_core/w[12] [29]),
	.I1(\top/processor/sha_core/w[13] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_138 )
);
defparam \top/processor/sha_core/n329_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s225  (
	.I0(\top/processor/sha_core/w[14] [29]),
	.I1(\top/processor/sha_core/w[15] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_139 )
);
defparam \top/processor/sha_core/n329_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s226  (
	.I0(\top/processor/sha_core/w[16] [29]),
	.I1(\top/processor/sha_core/w[17] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_140 )
);
defparam \top/processor/sha_core/n329_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s227  (
	.I0(\top/processor/sha_core/w[18] [29]),
	.I1(\top/processor/sha_core/w[19] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_141 )
);
defparam \top/processor/sha_core/n329_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s228  (
	.I0(\top/processor/sha_core/w[20] [29]),
	.I1(\top/processor/sha_core/w[21] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_142 )
);
defparam \top/processor/sha_core/n329_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s229  (
	.I0(\top/processor/sha_core/w[22] [29]),
	.I1(\top/processor/sha_core/w[23] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_143 )
);
defparam \top/processor/sha_core/n329_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s230  (
	.I0(\top/processor/sha_core/w[24] [29]),
	.I1(\top/processor/sha_core/w[25] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_144 )
);
defparam \top/processor/sha_core/n329_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s231  (
	.I0(\top/processor/sha_core/w[26] [29]),
	.I1(\top/processor/sha_core/w[27] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_145 )
);
defparam \top/processor/sha_core/n329_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s232  (
	.I0(\top/processor/sha_core/w[28] [29]),
	.I1(\top/processor/sha_core/w[29] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_146 )
);
defparam \top/processor/sha_core/n329_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s233  (
	.I0(\top/processor/sha_core/w[30] [29]),
	.I1(\top/processor/sha_core/w[31] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_147 )
);
defparam \top/processor/sha_core/n329_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s234  (
	.I0(\top/processor/sha_core/w[32] [29]),
	.I1(\top/processor/sha_core/w[33] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_148 )
);
defparam \top/processor/sha_core/n329_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s235  (
	.I0(\top/processor/sha_core/w[34] [29]),
	.I1(\top/processor/sha_core/w[35] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_149 )
);
defparam \top/processor/sha_core/n329_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s236  (
	.I0(\top/processor/sha_core/w[36] [29]),
	.I1(\top/processor/sha_core/w[37] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_150 )
);
defparam \top/processor/sha_core/n329_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s237  (
	.I0(\top/processor/sha_core/w[38] [29]),
	.I1(\top/processor/sha_core/w[39] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_151 )
);
defparam \top/processor/sha_core/n329_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s238  (
	.I0(\top/processor/sha_core/w[40] [29]),
	.I1(\top/processor/sha_core/w[41] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_152 )
);
defparam \top/processor/sha_core/n329_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s239  (
	.I0(\top/processor/sha_core/w[42] [29]),
	.I1(\top/processor/sha_core/w[43] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_153 )
);
defparam \top/processor/sha_core/n329_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s240  (
	.I0(\top/processor/sha_core/w[44] [29]),
	.I1(\top/processor/sha_core/w[45] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_154 )
);
defparam \top/processor/sha_core/n329_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s241  (
	.I0(\top/processor/sha_core/w[46] [29]),
	.I1(\top/processor/sha_core/w[47] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_155 )
);
defparam \top/processor/sha_core/n329_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s242  (
	.I0(\top/processor/sha_core/w[48] [29]),
	.I1(\top/processor/sha_core/w[49] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_156 )
);
defparam \top/processor/sha_core/n329_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s243  (
	.I0(\top/processor/sha_core/w[50] [29]),
	.I1(\top/processor/sha_core/w[51] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_157 )
);
defparam \top/processor/sha_core/n329_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s244  (
	.I0(\top/processor/sha_core/w[52] [29]),
	.I1(\top/processor/sha_core/w[53] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_158 )
);
defparam \top/processor/sha_core/n329_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s245  (
	.I0(\top/processor/sha_core/w[54] [29]),
	.I1(\top/processor/sha_core/w[55] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_159 )
);
defparam \top/processor/sha_core/n329_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s246  (
	.I0(\top/processor/sha_core/w[56] [29]),
	.I1(\top/processor/sha_core/w[57] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_160 )
);
defparam \top/processor/sha_core/n329_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s247  (
	.I0(\top/processor/sha_core/w[58] [29]),
	.I1(\top/processor/sha_core/w[59] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_161 )
);
defparam \top/processor/sha_core/n329_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s248  (
	.I0(\top/processor/sha_core/w[60] [29]),
	.I1(\top/processor/sha_core/w[61] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_162 )
);
defparam \top/processor/sha_core/n329_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s249  (
	.I0(\top/processor/sha_core/w[62] [29]),
	.I1(\top/processor/sha_core/w[63] [29]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n329_163 )
);
defparam \top/processor/sha_core/n329_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s218  (
	.I0(\top/processor/sha_core/w[0] [28]),
	.I1(\top/processor/sha_core/w[1] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_132 )
);
defparam \top/processor/sha_core/n330_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s219  (
	.I0(\top/processor/sha_core/w[2] [28]),
	.I1(\top/processor/sha_core/w[3] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_133 )
);
defparam \top/processor/sha_core/n330_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s220  (
	.I0(\top/processor/sha_core/w[4] [28]),
	.I1(\top/processor/sha_core/w[5] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_134 )
);
defparam \top/processor/sha_core/n330_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s221  (
	.I0(\top/processor/sha_core/w[6] [28]),
	.I1(\top/processor/sha_core/w[7] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_135 )
);
defparam \top/processor/sha_core/n330_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s222  (
	.I0(\top/processor/sha_core/w[8] [28]),
	.I1(\top/processor/sha_core/w[9] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_136 )
);
defparam \top/processor/sha_core/n330_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s223  (
	.I0(\top/processor/sha_core/w[10] [28]),
	.I1(\top/processor/sha_core/w[11] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_137 )
);
defparam \top/processor/sha_core/n330_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s224  (
	.I0(\top/processor/sha_core/w[12] [28]),
	.I1(\top/processor/sha_core/w[13] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_138 )
);
defparam \top/processor/sha_core/n330_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s225  (
	.I0(\top/processor/sha_core/w[14] [28]),
	.I1(\top/processor/sha_core/w[15] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_139 )
);
defparam \top/processor/sha_core/n330_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s226  (
	.I0(\top/processor/sha_core/w[16] [28]),
	.I1(\top/processor/sha_core/w[17] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_140 )
);
defparam \top/processor/sha_core/n330_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s227  (
	.I0(\top/processor/sha_core/w[18] [28]),
	.I1(\top/processor/sha_core/w[19] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_141 )
);
defparam \top/processor/sha_core/n330_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s228  (
	.I0(\top/processor/sha_core/w[20] [28]),
	.I1(\top/processor/sha_core/w[21] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_142 )
);
defparam \top/processor/sha_core/n330_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s229  (
	.I0(\top/processor/sha_core/w[22] [28]),
	.I1(\top/processor/sha_core/w[23] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_143 )
);
defparam \top/processor/sha_core/n330_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s230  (
	.I0(\top/processor/sha_core/w[24] [28]),
	.I1(\top/processor/sha_core/w[25] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_144 )
);
defparam \top/processor/sha_core/n330_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s231  (
	.I0(\top/processor/sha_core/w[26] [28]),
	.I1(\top/processor/sha_core/w[27] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_145 )
);
defparam \top/processor/sha_core/n330_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s232  (
	.I0(\top/processor/sha_core/w[28] [28]),
	.I1(\top/processor/sha_core/w[29] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_146 )
);
defparam \top/processor/sha_core/n330_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s233  (
	.I0(\top/processor/sha_core/w[30] [28]),
	.I1(\top/processor/sha_core/w[31] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_147 )
);
defparam \top/processor/sha_core/n330_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s234  (
	.I0(\top/processor/sha_core/w[32] [28]),
	.I1(\top/processor/sha_core/w[33] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_148 )
);
defparam \top/processor/sha_core/n330_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s235  (
	.I0(\top/processor/sha_core/w[34] [28]),
	.I1(\top/processor/sha_core/w[35] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_149 )
);
defparam \top/processor/sha_core/n330_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s236  (
	.I0(\top/processor/sha_core/w[36] [28]),
	.I1(\top/processor/sha_core/w[37] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_150 )
);
defparam \top/processor/sha_core/n330_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s237  (
	.I0(\top/processor/sha_core/w[38] [28]),
	.I1(\top/processor/sha_core/w[39] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_151 )
);
defparam \top/processor/sha_core/n330_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s238  (
	.I0(\top/processor/sha_core/w[40] [28]),
	.I1(\top/processor/sha_core/w[41] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_152 )
);
defparam \top/processor/sha_core/n330_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s239  (
	.I0(\top/processor/sha_core/w[42] [28]),
	.I1(\top/processor/sha_core/w[43] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_153 )
);
defparam \top/processor/sha_core/n330_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s240  (
	.I0(\top/processor/sha_core/w[44] [28]),
	.I1(\top/processor/sha_core/w[45] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_154 )
);
defparam \top/processor/sha_core/n330_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s241  (
	.I0(\top/processor/sha_core/w[46] [28]),
	.I1(\top/processor/sha_core/w[47] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_155 )
);
defparam \top/processor/sha_core/n330_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s242  (
	.I0(\top/processor/sha_core/w[48] [28]),
	.I1(\top/processor/sha_core/w[49] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_156 )
);
defparam \top/processor/sha_core/n330_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s243  (
	.I0(\top/processor/sha_core/w[50] [28]),
	.I1(\top/processor/sha_core/w[51] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_157 )
);
defparam \top/processor/sha_core/n330_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s244  (
	.I0(\top/processor/sha_core/w[52] [28]),
	.I1(\top/processor/sha_core/w[53] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_158 )
);
defparam \top/processor/sha_core/n330_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s245  (
	.I0(\top/processor/sha_core/w[54] [28]),
	.I1(\top/processor/sha_core/w[55] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_159 )
);
defparam \top/processor/sha_core/n330_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s246  (
	.I0(\top/processor/sha_core/w[56] [28]),
	.I1(\top/processor/sha_core/w[57] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_160 )
);
defparam \top/processor/sha_core/n330_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s247  (
	.I0(\top/processor/sha_core/w[58] [28]),
	.I1(\top/processor/sha_core/w[59] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_161 )
);
defparam \top/processor/sha_core/n330_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s248  (
	.I0(\top/processor/sha_core/w[60] [28]),
	.I1(\top/processor/sha_core/w[61] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_162 )
);
defparam \top/processor/sha_core/n330_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s249  (
	.I0(\top/processor/sha_core/w[62] [28]),
	.I1(\top/processor/sha_core/w[63] [28]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n330_163 )
);
defparam \top/processor/sha_core/n330_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s218  (
	.I0(\top/processor/sha_core/w[0] [27]),
	.I1(\top/processor/sha_core/w[1] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_132 )
);
defparam \top/processor/sha_core/n331_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s219  (
	.I0(\top/processor/sha_core/w[2] [27]),
	.I1(\top/processor/sha_core/w[3] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_133 )
);
defparam \top/processor/sha_core/n331_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s220  (
	.I0(\top/processor/sha_core/w[4] [27]),
	.I1(\top/processor/sha_core/w[5] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_134 )
);
defparam \top/processor/sha_core/n331_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s221  (
	.I0(\top/processor/sha_core/w[6] [27]),
	.I1(\top/processor/sha_core/w[7] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_135 )
);
defparam \top/processor/sha_core/n331_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s222  (
	.I0(\top/processor/sha_core/w[8] [27]),
	.I1(\top/processor/sha_core/w[9] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_136 )
);
defparam \top/processor/sha_core/n331_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s223  (
	.I0(\top/processor/sha_core/w[10] [27]),
	.I1(\top/processor/sha_core/w[11] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_137 )
);
defparam \top/processor/sha_core/n331_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s224  (
	.I0(\top/processor/sha_core/w[12] [27]),
	.I1(\top/processor/sha_core/w[13] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_138 )
);
defparam \top/processor/sha_core/n331_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s225  (
	.I0(\top/processor/sha_core/w[14] [27]),
	.I1(\top/processor/sha_core/w[15] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_139 )
);
defparam \top/processor/sha_core/n331_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s226  (
	.I0(\top/processor/sha_core/w[16] [27]),
	.I1(\top/processor/sha_core/w[17] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_140 )
);
defparam \top/processor/sha_core/n331_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s227  (
	.I0(\top/processor/sha_core/w[18] [27]),
	.I1(\top/processor/sha_core/w[19] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_141 )
);
defparam \top/processor/sha_core/n331_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s228  (
	.I0(\top/processor/sha_core/w[20] [27]),
	.I1(\top/processor/sha_core/w[21] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_142 )
);
defparam \top/processor/sha_core/n331_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s229  (
	.I0(\top/processor/sha_core/w[22] [27]),
	.I1(\top/processor/sha_core/w[23] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_143 )
);
defparam \top/processor/sha_core/n331_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s230  (
	.I0(\top/processor/sha_core/w[24] [27]),
	.I1(\top/processor/sha_core/w[25] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_144 )
);
defparam \top/processor/sha_core/n331_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s231  (
	.I0(\top/processor/sha_core/w[26] [27]),
	.I1(\top/processor/sha_core/w[27] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_145 )
);
defparam \top/processor/sha_core/n331_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s232  (
	.I0(\top/processor/sha_core/w[28] [27]),
	.I1(\top/processor/sha_core/w[29] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_146 )
);
defparam \top/processor/sha_core/n331_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s233  (
	.I0(\top/processor/sha_core/w[30] [27]),
	.I1(\top/processor/sha_core/w[31] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_147 )
);
defparam \top/processor/sha_core/n331_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s234  (
	.I0(\top/processor/sha_core/w[32] [27]),
	.I1(\top/processor/sha_core/w[33] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_148 )
);
defparam \top/processor/sha_core/n331_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s235  (
	.I0(\top/processor/sha_core/w[34] [27]),
	.I1(\top/processor/sha_core/w[35] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_149 )
);
defparam \top/processor/sha_core/n331_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s236  (
	.I0(\top/processor/sha_core/w[36] [27]),
	.I1(\top/processor/sha_core/w[37] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_150 )
);
defparam \top/processor/sha_core/n331_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s237  (
	.I0(\top/processor/sha_core/w[38] [27]),
	.I1(\top/processor/sha_core/w[39] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_151 )
);
defparam \top/processor/sha_core/n331_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s238  (
	.I0(\top/processor/sha_core/w[40] [27]),
	.I1(\top/processor/sha_core/w[41] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_152 )
);
defparam \top/processor/sha_core/n331_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s239  (
	.I0(\top/processor/sha_core/w[42] [27]),
	.I1(\top/processor/sha_core/w[43] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_153 )
);
defparam \top/processor/sha_core/n331_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s240  (
	.I0(\top/processor/sha_core/w[44] [27]),
	.I1(\top/processor/sha_core/w[45] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_154 )
);
defparam \top/processor/sha_core/n331_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s241  (
	.I0(\top/processor/sha_core/w[46] [27]),
	.I1(\top/processor/sha_core/w[47] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_155 )
);
defparam \top/processor/sha_core/n331_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s242  (
	.I0(\top/processor/sha_core/w[48] [27]),
	.I1(\top/processor/sha_core/w[49] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_156 )
);
defparam \top/processor/sha_core/n331_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s243  (
	.I0(\top/processor/sha_core/w[50] [27]),
	.I1(\top/processor/sha_core/w[51] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_157 )
);
defparam \top/processor/sha_core/n331_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s244  (
	.I0(\top/processor/sha_core/w[52] [27]),
	.I1(\top/processor/sha_core/w[53] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_158 )
);
defparam \top/processor/sha_core/n331_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s245  (
	.I0(\top/processor/sha_core/w[54] [27]),
	.I1(\top/processor/sha_core/w[55] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_159 )
);
defparam \top/processor/sha_core/n331_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s246  (
	.I0(\top/processor/sha_core/w[56] [27]),
	.I1(\top/processor/sha_core/w[57] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_160 )
);
defparam \top/processor/sha_core/n331_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s247  (
	.I0(\top/processor/sha_core/w[58] [27]),
	.I1(\top/processor/sha_core/w[59] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_161 )
);
defparam \top/processor/sha_core/n331_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s248  (
	.I0(\top/processor/sha_core/w[60] [27]),
	.I1(\top/processor/sha_core/w[61] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_162 )
);
defparam \top/processor/sha_core/n331_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s249  (
	.I0(\top/processor/sha_core/w[62] [27]),
	.I1(\top/processor/sha_core/w[63] [27]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n331_163 )
);
defparam \top/processor/sha_core/n331_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s218  (
	.I0(\top/processor/sha_core/w[0] [26]),
	.I1(\top/processor/sha_core/w[1] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_132 )
);
defparam \top/processor/sha_core/n332_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s219  (
	.I0(\top/processor/sha_core/w[2] [26]),
	.I1(\top/processor/sha_core/w[3] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_133 )
);
defparam \top/processor/sha_core/n332_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s220  (
	.I0(\top/processor/sha_core/w[4] [26]),
	.I1(\top/processor/sha_core/w[5] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_134 )
);
defparam \top/processor/sha_core/n332_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s221  (
	.I0(\top/processor/sha_core/w[6] [26]),
	.I1(\top/processor/sha_core/w[7] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_135 )
);
defparam \top/processor/sha_core/n332_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s222  (
	.I0(\top/processor/sha_core/w[8] [26]),
	.I1(\top/processor/sha_core/w[9] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_136 )
);
defparam \top/processor/sha_core/n332_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s223  (
	.I0(\top/processor/sha_core/w[10] [26]),
	.I1(\top/processor/sha_core/w[11] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_137 )
);
defparam \top/processor/sha_core/n332_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s224  (
	.I0(\top/processor/sha_core/w[12] [26]),
	.I1(\top/processor/sha_core/w[13] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_138 )
);
defparam \top/processor/sha_core/n332_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s225  (
	.I0(\top/processor/sha_core/w[14] [26]),
	.I1(\top/processor/sha_core/w[15] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_139 )
);
defparam \top/processor/sha_core/n332_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s226  (
	.I0(\top/processor/sha_core/w[16] [26]),
	.I1(\top/processor/sha_core/w[17] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_140 )
);
defparam \top/processor/sha_core/n332_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s227  (
	.I0(\top/processor/sha_core/w[18] [26]),
	.I1(\top/processor/sha_core/w[19] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_141 )
);
defparam \top/processor/sha_core/n332_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s228  (
	.I0(\top/processor/sha_core/w[20] [26]),
	.I1(\top/processor/sha_core/w[21] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_142 )
);
defparam \top/processor/sha_core/n332_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s229  (
	.I0(\top/processor/sha_core/w[22] [26]),
	.I1(\top/processor/sha_core/w[23] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_143 )
);
defparam \top/processor/sha_core/n332_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s230  (
	.I0(\top/processor/sha_core/w[24] [26]),
	.I1(\top/processor/sha_core/w[25] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_144 )
);
defparam \top/processor/sha_core/n332_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s231  (
	.I0(\top/processor/sha_core/w[26] [26]),
	.I1(\top/processor/sha_core/w[27] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_145 )
);
defparam \top/processor/sha_core/n332_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s232  (
	.I0(\top/processor/sha_core/w[28] [26]),
	.I1(\top/processor/sha_core/w[29] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_146 )
);
defparam \top/processor/sha_core/n332_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s233  (
	.I0(\top/processor/sha_core/w[30] [26]),
	.I1(\top/processor/sha_core/w[31] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_147 )
);
defparam \top/processor/sha_core/n332_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s234  (
	.I0(\top/processor/sha_core/w[32] [26]),
	.I1(\top/processor/sha_core/w[33] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_148 )
);
defparam \top/processor/sha_core/n332_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s235  (
	.I0(\top/processor/sha_core/w[34] [26]),
	.I1(\top/processor/sha_core/w[35] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_149 )
);
defparam \top/processor/sha_core/n332_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s236  (
	.I0(\top/processor/sha_core/w[36] [26]),
	.I1(\top/processor/sha_core/w[37] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_150 )
);
defparam \top/processor/sha_core/n332_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s237  (
	.I0(\top/processor/sha_core/w[38] [26]),
	.I1(\top/processor/sha_core/w[39] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_151 )
);
defparam \top/processor/sha_core/n332_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s238  (
	.I0(\top/processor/sha_core/w[40] [26]),
	.I1(\top/processor/sha_core/w[41] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_152 )
);
defparam \top/processor/sha_core/n332_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s239  (
	.I0(\top/processor/sha_core/w[42] [26]),
	.I1(\top/processor/sha_core/w[43] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_153 )
);
defparam \top/processor/sha_core/n332_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s240  (
	.I0(\top/processor/sha_core/w[44] [26]),
	.I1(\top/processor/sha_core/w[45] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_154 )
);
defparam \top/processor/sha_core/n332_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s241  (
	.I0(\top/processor/sha_core/w[46] [26]),
	.I1(\top/processor/sha_core/w[47] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_155 )
);
defparam \top/processor/sha_core/n332_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s242  (
	.I0(\top/processor/sha_core/w[48] [26]),
	.I1(\top/processor/sha_core/w[49] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_156 )
);
defparam \top/processor/sha_core/n332_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s243  (
	.I0(\top/processor/sha_core/w[50] [26]),
	.I1(\top/processor/sha_core/w[51] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_157 )
);
defparam \top/processor/sha_core/n332_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s244  (
	.I0(\top/processor/sha_core/w[52] [26]),
	.I1(\top/processor/sha_core/w[53] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_158 )
);
defparam \top/processor/sha_core/n332_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s245  (
	.I0(\top/processor/sha_core/w[54] [26]),
	.I1(\top/processor/sha_core/w[55] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_159 )
);
defparam \top/processor/sha_core/n332_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s246  (
	.I0(\top/processor/sha_core/w[56] [26]),
	.I1(\top/processor/sha_core/w[57] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_160 )
);
defparam \top/processor/sha_core/n332_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s247  (
	.I0(\top/processor/sha_core/w[58] [26]),
	.I1(\top/processor/sha_core/w[59] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_161 )
);
defparam \top/processor/sha_core/n332_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s248  (
	.I0(\top/processor/sha_core/w[60] [26]),
	.I1(\top/processor/sha_core/w[61] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_162 )
);
defparam \top/processor/sha_core/n332_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s249  (
	.I0(\top/processor/sha_core/w[62] [26]),
	.I1(\top/processor/sha_core/w[63] [26]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n332_163 )
);
defparam \top/processor/sha_core/n332_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s218  (
	.I0(\top/processor/sha_core/w[0] [25]),
	.I1(\top/processor/sha_core/w[1] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_132 )
);
defparam \top/processor/sha_core/n333_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s219  (
	.I0(\top/processor/sha_core/w[2] [25]),
	.I1(\top/processor/sha_core/w[3] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_133 )
);
defparam \top/processor/sha_core/n333_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s220  (
	.I0(\top/processor/sha_core/w[4] [25]),
	.I1(\top/processor/sha_core/w[5] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_134 )
);
defparam \top/processor/sha_core/n333_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s221  (
	.I0(\top/processor/sha_core/w[6] [25]),
	.I1(\top/processor/sha_core/w[7] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_135 )
);
defparam \top/processor/sha_core/n333_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s222  (
	.I0(\top/processor/sha_core/w[8] [25]),
	.I1(\top/processor/sha_core/w[9] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_136 )
);
defparam \top/processor/sha_core/n333_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s223  (
	.I0(\top/processor/sha_core/w[10] [25]),
	.I1(\top/processor/sha_core/w[11] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_137 )
);
defparam \top/processor/sha_core/n333_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s224  (
	.I0(\top/processor/sha_core/w[12] [25]),
	.I1(\top/processor/sha_core/w[13] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_138 )
);
defparam \top/processor/sha_core/n333_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s225  (
	.I0(\top/processor/sha_core/w[14] [25]),
	.I1(\top/processor/sha_core/w[15] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_139 )
);
defparam \top/processor/sha_core/n333_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s226  (
	.I0(\top/processor/sha_core/w[16] [25]),
	.I1(\top/processor/sha_core/w[17] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_140 )
);
defparam \top/processor/sha_core/n333_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s227  (
	.I0(\top/processor/sha_core/w[18] [25]),
	.I1(\top/processor/sha_core/w[19] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_141 )
);
defparam \top/processor/sha_core/n333_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s228  (
	.I0(\top/processor/sha_core/w[20] [25]),
	.I1(\top/processor/sha_core/w[21] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_142 )
);
defparam \top/processor/sha_core/n333_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s229  (
	.I0(\top/processor/sha_core/w[22] [25]),
	.I1(\top/processor/sha_core/w[23] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_143 )
);
defparam \top/processor/sha_core/n333_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s230  (
	.I0(\top/processor/sha_core/w[24] [25]),
	.I1(\top/processor/sha_core/w[25] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_144 )
);
defparam \top/processor/sha_core/n333_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s231  (
	.I0(\top/processor/sha_core/w[26] [25]),
	.I1(\top/processor/sha_core/w[27] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_145 )
);
defparam \top/processor/sha_core/n333_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s232  (
	.I0(\top/processor/sha_core/w[28] [25]),
	.I1(\top/processor/sha_core/w[29] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_146 )
);
defparam \top/processor/sha_core/n333_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s233  (
	.I0(\top/processor/sha_core/w[30] [25]),
	.I1(\top/processor/sha_core/w[31] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_147 )
);
defparam \top/processor/sha_core/n333_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s234  (
	.I0(\top/processor/sha_core/w[32] [25]),
	.I1(\top/processor/sha_core/w[33] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_148 )
);
defparam \top/processor/sha_core/n333_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s235  (
	.I0(\top/processor/sha_core/w[34] [25]),
	.I1(\top/processor/sha_core/w[35] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_149 )
);
defparam \top/processor/sha_core/n333_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s236  (
	.I0(\top/processor/sha_core/w[36] [25]),
	.I1(\top/processor/sha_core/w[37] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_150 )
);
defparam \top/processor/sha_core/n333_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s237  (
	.I0(\top/processor/sha_core/w[38] [25]),
	.I1(\top/processor/sha_core/w[39] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_151 )
);
defparam \top/processor/sha_core/n333_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s238  (
	.I0(\top/processor/sha_core/w[40] [25]),
	.I1(\top/processor/sha_core/w[41] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_152 )
);
defparam \top/processor/sha_core/n333_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s239  (
	.I0(\top/processor/sha_core/w[42] [25]),
	.I1(\top/processor/sha_core/w[43] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_153 )
);
defparam \top/processor/sha_core/n333_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s240  (
	.I0(\top/processor/sha_core/w[44] [25]),
	.I1(\top/processor/sha_core/w[45] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_154 )
);
defparam \top/processor/sha_core/n333_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s241  (
	.I0(\top/processor/sha_core/w[46] [25]),
	.I1(\top/processor/sha_core/w[47] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_155 )
);
defparam \top/processor/sha_core/n333_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s242  (
	.I0(\top/processor/sha_core/w[48] [25]),
	.I1(\top/processor/sha_core/w[49] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_156 )
);
defparam \top/processor/sha_core/n333_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s243  (
	.I0(\top/processor/sha_core/w[50] [25]),
	.I1(\top/processor/sha_core/w[51] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_157 )
);
defparam \top/processor/sha_core/n333_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s244  (
	.I0(\top/processor/sha_core/w[52] [25]),
	.I1(\top/processor/sha_core/w[53] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_158 )
);
defparam \top/processor/sha_core/n333_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s245  (
	.I0(\top/processor/sha_core/w[54] [25]),
	.I1(\top/processor/sha_core/w[55] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_159 )
);
defparam \top/processor/sha_core/n333_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s246  (
	.I0(\top/processor/sha_core/w[56] [25]),
	.I1(\top/processor/sha_core/w[57] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_160 )
);
defparam \top/processor/sha_core/n333_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s247  (
	.I0(\top/processor/sha_core/w[58] [25]),
	.I1(\top/processor/sha_core/w[59] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_161 )
);
defparam \top/processor/sha_core/n333_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s248  (
	.I0(\top/processor/sha_core/w[60] [25]),
	.I1(\top/processor/sha_core/w[61] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_162 )
);
defparam \top/processor/sha_core/n333_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s249  (
	.I0(\top/processor/sha_core/w[62] [25]),
	.I1(\top/processor/sha_core/w[63] [25]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n333_163 )
);
defparam \top/processor/sha_core/n333_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s218  (
	.I0(\top/processor/sha_core/w[0] [24]),
	.I1(\top/processor/sha_core/w[1] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_132 )
);
defparam \top/processor/sha_core/n334_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s219  (
	.I0(\top/processor/sha_core/w[2] [24]),
	.I1(\top/processor/sha_core/w[3] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_133 )
);
defparam \top/processor/sha_core/n334_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s220  (
	.I0(\top/processor/sha_core/w[4] [24]),
	.I1(\top/processor/sha_core/w[5] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_134 )
);
defparam \top/processor/sha_core/n334_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s221  (
	.I0(\top/processor/sha_core/w[6] [24]),
	.I1(\top/processor/sha_core/w[7] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_135 )
);
defparam \top/processor/sha_core/n334_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s222  (
	.I0(\top/processor/sha_core/w[8] [24]),
	.I1(\top/processor/sha_core/w[9] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_136 )
);
defparam \top/processor/sha_core/n334_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s223  (
	.I0(\top/processor/sha_core/w[10] [24]),
	.I1(\top/processor/sha_core/w[11] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_137 )
);
defparam \top/processor/sha_core/n334_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s224  (
	.I0(\top/processor/sha_core/w[12] [24]),
	.I1(\top/processor/sha_core/w[13] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_138 )
);
defparam \top/processor/sha_core/n334_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s225  (
	.I0(\top/processor/sha_core/w[14] [24]),
	.I1(\top/processor/sha_core/w[15] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_139 )
);
defparam \top/processor/sha_core/n334_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s226  (
	.I0(\top/processor/sha_core/w[16] [24]),
	.I1(\top/processor/sha_core/w[17] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_140 )
);
defparam \top/processor/sha_core/n334_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s227  (
	.I0(\top/processor/sha_core/w[18] [24]),
	.I1(\top/processor/sha_core/w[19] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_141 )
);
defparam \top/processor/sha_core/n334_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s228  (
	.I0(\top/processor/sha_core/w[20] [24]),
	.I1(\top/processor/sha_core/w[21] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_142 )
);
defparam \top/processor/sha_core/n334_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s229  (
	.I0(\top/processor/sha_core/w[22] [24]),
	.I1(\top/processor/sha_core/w[23] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_143 )
);
defparam \top/processor/sha_core/n334_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s230  (
	.I0(\top/processor/sha_core/w[24] [24]),
	.I1(\top/processor/sha_core/w[25] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_144 )
);
defparam \top/processor/sha_core/n334_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s231  (
	.I0(\top/processor/sha_core/w[26] [24]),
	.I1(\top/processor/sha_core/w[27] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_145 )
);
defparam \top/processor/sha_core/n334_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s232  (
	.I0(\top/processor/sha_core/w[28] [24]),
	.I1(\top/processor/sha_core/w[29] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_146 )
);
defparam \top/processor/sha_core/n334_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s233  (
	.I0(\top/processor/sha_core/w[30] [24]),
	.I1(\top/processor/sha_core/w[31] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_147 )
);
defparam \top/processor/sha_core/n334_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s234  (
	.I0(\top/processor/sha_core/w[32] [24]),
	.I1(\top/processor/sha_core/w[33] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_148 )
);
defparam \top/processor/sha_core/n334_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s235  (
	.I0(\top/processor/sha_core/w[34] [24]),
	.I1(\top/processor/sha_core/w[35] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_149 )
);
defparam \top/processor/sha_core/n334_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s236  (
	.I0(\top/processor/sha_core/w[36] [24]),
	.I1(\top/processor/sha_core/w[37] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_150 )
);
defparam \top/processor/sha_core/n334_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s237  (
	.I0(\top/processor/sha_core/w[38] [24]),
	.I1(\top/processor/sha_core/w[39] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_151 )
);
defparam \top/processor/sha_core/n334_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s238  (
	.I0(\top/processor/sha_core/w[40] [24]),
	.I1(\top/processor/sha_core/w[41] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_152 )
);
defparam \top/processor/sha_core/n334_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s239  (
	.I0(\top/processor/sha_core/w[42] [24]),
	.I1(\top/processor/sha_core/w[43] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_153 )
);
defparam \top/processor/sha_core/n334_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s240  (
	.I0(\top/processor/sha_core/w[44] [24]),
	.I1(\top/processor/sha_core/w[45] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_154 )
);
defparam \top/processor/sha_core/n334_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s241  (
	.I0(\top/processor/sha_core/w[46] [24]),
	.I1(\top/processor/sha_core/w[47] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_155 )
);
defparam \top/processor/sha_core/n334_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s242  (
	.I0(\top/processor/sha_core/w[48] [24]),
	.I1(\top/processor/sha_core/w[49] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_156 )
);
defparam \top/processor/sha_core/n334_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s243  (
	.I0(\top/processor/sha_core/w[50] [24]),
	.I1(\top/processor/sha_core/w[51] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_157 )
);
defparam \top/processor/sha_core/n334_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s244  (
	.I0(\top/processor/sha_core/w[52] [24]),
	.I1(\top/processor/sha_core/w[53] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_158 )
);
defparam \top/processor/sha_core/n334_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s245  (
	.I0(\top/processor/sha_core/w[54] [24]),
	.I1(\top/processor/sha_core/w[55] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_159 )
);
defparam \top/processor/sha_core/n334_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s246  (
	.I0(\top/processor/sha_core/w[56] [24]),
	.I1(\top/processor/sha_core/w[57] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_160 )
);
defparam \top/processor/sha_core/n334_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s247  (
	.I0(\top/processor/sha_core/w[58] [24]),
	.I1(\top/processor/sha_core/w[59] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_161 )
);
defparam \top/processor/sha_core/n334_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s248  (
	.I0(\top/processor/sha_core/w[60] [24]),
	.I1(\top/processor/sha_core/w[61] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_162 )
);
defparam \top/processor/sha_core/n334_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s249  (
	.I0(\top/processor/sha_core/w[62] [24]),
	.I1(\top/processor/sha_core/w[63] [24]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n334_163 )
);
defparam \top/processor/sha_core/n334_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s218  (
	.I0(\top/processor/sha_core/w[0] [23]),
	.I1(\top/processor/sha_core/w[1] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_132 )
);
defparam \top/processor/sha_core/n335_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s219  (
	.I0(\top/processor/sha_core/w[2] [23]),
	.I1(\top/processor/sha_core/w[3] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_133 )
);
defparam \top/processor/sha_core/n335_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s220  (
	.I0(\top/processor/sha_core/w[4] [23]),
	.I1(\top/processor/sha_core/w[5] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_134 )
);
defparam \top/processor/sha_core/n335_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s221  (
	.I0(\top/processor/sha_core/w[6] [23]),
	.I1(\top/processor/sha_core/w[7] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_135 )
);
defparam \top/processor/sha_core/n335_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s222  (
	.I0(\top/processor/sha_core/w[8] [23]),
	.I1(\top/processor/sha_core/w[9] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_136 )
);
defparam \top/processor/sha_core/n335_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s223  (
	.I0(\top/processor/sha_core/w[10] [23]),
	.I1(\top/processor/sha_core/w[11] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_137 )
);
defparam \top/processor/sha_core/n335_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s224  (
	.I0(\top/processor/sha_core/w[12] [23]),
	.I1(\top/processor/sha_core/w[13] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_138 )
);
defparam \top/processor/sha_core/n335_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s225  (
	.I0(\top/processor/sha_core/w[14] [23]),
	.I1(\top/processor/sha_core/w[15] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_139 )
);
defparam \top/processor/sha_core/n335_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s226  (
	.I0(\top/processor/sha_core/w[16] [23]),
	.I1(\top/processor/sha_core/w[17] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_140 )
);
defparam \top/processor/sha_core/n335_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s227  (
	.I0(\top/processor/sha_core/w[18] [23]),
	.I1(\top/processor/sha_core/w[19] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_141 )
);
defparam \top/processor/sha_core/n335_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s228  (
	.I0(\top/processor/sha_core/w[20] [23]),
	.I1(\top/processor/sha_core/w[21] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_142 )
);
defparam \top/processor/sha_core/n335_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s229  (
	.I0(\top/processor/sha_core/w[22] [23]),
	.I1(\top/processor/sha_core/w[23] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_143 )
);
defparam \top/processor/sha_core/n335_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s230  (
	.I0(\top/processor/sha_core/w[24] [23]),
	.I1(\top/processor/sha_core/w[25] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_144 )
);
defparam \top/processor/sha_core/n335_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s231  (
	.I0(\top/processor/sha_core/w[26] [23]),
	.I1(\top/processor/sha_core/w[27] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_145 )
);
defparam \top/processor/sha_core/n335_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s232  (
	.I0(\top/processor/sha_core/w[28] [23]),
	.I1(\top/processor/sha_core/w[29] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_146 )
);
defparam \top/processor/sha_core/n335_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s233  (
	.I0(\top/processor/sha_core/w[30] [23]),
	.I1(\top/processor/sha_core/w[31] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_147 )
);
defparam \top/processor/sha_core/n335_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s234  (
	.I0(\top/processor/sha_core/w[32] [23]),
	.I1(\top/processor/sha_core/w[33] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_148 )
);
defparam \top/processor/sha_core/n335_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s235  (
	.I0(\top/processor/sha_core/w[34] [23]),
	.I1(\top/processor/sha_core/w[35] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_149 )
);
defparam \top/processor/sha_core/n335_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s236  (
	.I0(\top/processor/sha_core/w[36] [23]),
	.I1(\top/processor/sha_core/w[37] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_150 )
);
defparam \top/processor/sha_core/n335_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s237  (
	.I0(\top/processor/sha_core/w[38] [23]),
	.I1(\top/processor/sha_core/w[39] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_151 )
);
defparam \top/processor/sha_core/n335_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s238  (
	.I0(\top/processor/sha_core/w[40] [23]),
	.I1(\top/processor/sha_core/w[41] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_152 )
);
defparam \top/processor/sha_core/n335_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s239  (
	.I0(\top/processor/sha_core/w[42] [23]),
	.I1(\top/processor/sha_core/w[43] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_153 )
);
defparam \top/processor/sha_core/n335_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s240  (
	.I0(\top/processor/sha_core/w[44] [23]),
	.I1(\top/processor/sha_core/w[45] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_154 )
);
defparam \top/processor/sha_core/n335_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s241  (
	.I0(\top/processor/sha_core/w[46] [23]),
	.I1(\top/processor/sha_core/w[47] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_155 )
);
defparam \top/processor/sha_core/n335_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s242  (
	.I0(\top/processor/sha_core/w[48] [23]),
	.I1(\top/processor/sha_core/w[49] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_156 )
);
defparam \top/processor/sha_core/n335_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s243  (
	.I0(\top/processor/sha_core/w[50] [23]),
	.I1(\top/processor/sha_core/w[51] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_157 )
);
defparam \top/processor/sha_core/n335_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s244  (
	.I0(\top/processor/sha_core/w[52] [23]),
	.I1(\top/processor/sha_core/w[53] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_158 )
);
defparam \top/processor/sha_core/n335_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s245  (
	.I0(\top/processor/sha_core/w[54] [23]),
	.I1(\top/processor/sha_core/w[55] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_159 )
);
defparam \top/processor/sha_core/n335_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s246  (
	.I0(\top/processor/sha_core/w[56] [23]),
	.I1(\top/processor/sha_core/w[57] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_160 )
);
defparam \top/processor/sha_core/n335_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s247  (
	.I0(\top/processor/sha_core/w[58] [23]),
	.I1(\top/processor/sha_core/w[59] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_161 )
);
defparam \top/processor/sha_core/n335_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s248  (
	.I0(\top/processor/sha_core/w[60] [23]),
	.I1(\top/processor/sha_core/w[61] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_162 )
);
defparam \top/processor/sha_core/n335_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s249  (
	.I0(\top/processor/sha_core/w[62] [23]),
	.I1(\top/processor/sha_core/w[63] [23]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n335_163 )
);
defparam \top/processor/sha_core/n335_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s218  (
	.I0(\top/processor/sha_core/w[0] [22]),
	.I1(\top/processor/sha_core/w[1] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_132 )
);
defparam \top/processor/sha_core/n336_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s219  (
	.I0(\top/processor/sha_core/w[2] [22]),
	.I1(\top/processor/sha_core/w[3] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_133 )
);
defparam \top/processor/sha_core/n336_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s220  (
	.I0(\top/processor/sha_core/w[4] [22]),
	.I1(\top/processor/sha_core/w[5] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_134 )
);
defparam \top/processor/sha_core/n336_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s221  (
	.I0(\top/processor/sha_core/w[6] [22]),
	.I1(\top/processor/sha_core/w[7] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_135 )
);
defparam \top/processor/sha_core/n336_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s222  (
	.I0(\top/processor/sha_core/w[8] [22]),
	.I1(\top/processor/sha_core/w[9] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_136 )
);
defparam \top/processor/sha_core/n336_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s223  (
	.I0(\top/processor/sha_core/w[10] [22]),
	.I1(\top/processor/sha_core/w[11] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_137 )
);
defparam \top/processor/sha_core/n336_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s224  (
	.I0(\top/processor/sha_core/w[12] [22]),
	.I1(\top/processor/sha_core/w[13] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_138 )
);
defparam \top/processor/sha_core/n336_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s225  (
	.I0(\top/processor/sha_core/w[14] [22]),
	.I1(\top/processor/sha_core/w[15] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_139 )
);
defparam \top/processor/sha_core/n336_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s226  (
	.I0(\top/processor/sha_core/w[16] [22]),
	.I1(\top/processor/sha_core/w[17] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_140 )
);
defparam \top/processor/sha_core/n336_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s227  (
	.I0(\top/processor/sha_core/w[18] [22]),
	.I1(\top/processor/sha_core/w[19] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_141 )
);
defparam \top/processor/sha_core/n336_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s228  (
	.I0(\top/processor/sha_core/w[20] [22]),
	.I1(\top/processor/sha_core/w[21] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_142 )
);
defparam \top/processor/sha_core/n336_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s229  (
	.I0(\top/processor/sha_core/w[22] [22]),
	.I1(\top/processor/sha_core/w[23] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_143 )
);
defparam \top/processor/sha_core/n336_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s230  (
	.I0(\top/processor/sha_core/w[24] [22]),
	.I1(\top/processor/sha_core/w[25] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_144 )
);
defparam \top/processor/sha_core/n336_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s231  (
	.I0(\top/processor/sha_core/w[26] [22]),
	.I1(\top/processor/sha_core/w[27] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_145 )
);
defparam \top/processor/sha_core/n336_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s232  (
	.I0(\top/processor/sha_core/w[28] [22]),
	.I1(\top/processor/sha_core/w[29] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_146 )
);
defparam \top/processor/sha_core/n336_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s233  (
	.I0(\top/processor/sha_core/w[30] [22]),
	.I1(\top/processor/sha_core/w[31] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_147 )
);
defparam \top/processor/sha_core/n336_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s234  (
	.I0(\top/processor/sha_core/w[32] [22]),
	.I1(\top/processor/sha_core/w[33] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_148 )
);
defparam \top/processor/sha_core/n336_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s235  (
	.I0(\top/processor/sha_core/w[34] [22]),
	.I1(\top/processor/sha_core/w[35] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_149 )
);
defparam \top/processor/sha_core/n336_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s236  (
	.I0(\top/processor/sha_core/w[36] [22]),
	.I1(\top/processor/sha_core/w[37] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_150 )
);
defparam \top/processor/sha_core/n336_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s237  (
	.I0(\top/processor/sha_core/w[38] [22]),
	.I1(\top/processor/sha_core/w[39] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_151 )
);
defparam \top/processor/sha_core/n336_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s238  (
	.I0(\top/processor/sha_core/w[40] [22]),
	.I1(\top/processor/sha_core/w[41] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_152 )
);
defparam \top/processor/sha_core/n336_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s239  (
	.I0(\top/processor/sha_core/w[42] [22]),
	.I1(\top/processor/sha_core/w[43] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_153 )
);
defparam \top/processor/sha_core/n336_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s240  (
	.I0(\top/processor/sha_core/w[44] [22]),
	.I1(\top/processor/sha_core/w[45] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_154 )
);
defparam \top/processor/sha_core/n336_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s241  (
	.I0(\top/processor/sha_core/w[46] [22]),
	.I1(\top/processor/sha_core/w[47] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_155 )
);
defparam \top/processor/sha_core/n336_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s242  (
	.I0(\top/processor/sha_core/w[48] [22]),
	.I1(\top/processor/sha_core/w[49] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_156 )
);
defparam \top/processor/sha_core/n336_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s243  (
	.I0(\top/processor/sha_core/w[50] [22]),
	.I1(\top/processor/sha_core/w[51] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_157 )
);
defparam \top/processor/sha_core/n336_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s244  (
	.I0(\top/processor/sha_core/w[52] [22]),
	.I1(\top/processor/sha_core/w[53] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_158 )
);
defparam \top/processor/sha_core/n336_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s245  (
	.I0(\top/processor/sha_core/w[54] [22]),
	.I1(\top/processor/sha_core/w[55] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_159 )
);
defparam \top/processor/sha_core/n336_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s246  (
	.I0(\top/processor/sha_core/w[56] [22]),
	.I1(\top/processor/sha_core/w[57] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_160 )
);
defparam \top/processor/sha_core/n336_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s247  (
	.I0(\top/processor/sha_core/w[58] [22]),
	.I1(\top/processor/sha_core/w[59] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_161 )
);
defparam \top/processor/sha_core/n336_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s248  (
	.I0(\top/processor/sha_core/w[60] [22]),
	.I1(\top/processor/sha_core/w[61] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_162 )
);
defparam \top/processor/sha_core/n336_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s249  (
	.I0(\top/processor/sha_core/w[62] [22]),
	.I1(\top/processor/sha_core/w[63] [22]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n336_163 )
);
defparam \top/processor/sha_core/n336_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s218  (
	.I0(\top/processor/sha_core/w[0] [21]),
	.I1(\top/processor/sha_core/w[1] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_132 )
);
defparam \top/processor/sha_core/n337_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s219  (
	.I0(\top/processor/sha_core/w[2] [21]),
	.I1(\top/processor/sha_core/w[3] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_133 )
);
defparam \top/processor/sha_core/n337_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s220  (
	.I0(\top/processor/sha_core/w[4] [21]),
	.I1(\top/processor/sha_core/w[5] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_134 )
);
defparam \top/processor/sha_core/n337_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s221  (
	.I0(\top/processor/sha_core/w[6] [21]),
	.I1(\top/processor/sha_core/w[7] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_135 )
);
defparam \top/processor/sha_core/n337_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s222  (
	.I0(\top/processor/sha_core/w[8] [21]),
	.I1(\top/processor/sha_core/w[9] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_136 )
);
defparam \top/processor/sha_core/n337_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s223  (
	.I0(\top/processor/sha_core/w[10] [21]),
	.I1(\top/processor/sha_core/w[11] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_137 )
);
defparam \top/processor/sha_core/n337_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s224  (
	.I0(\top/processor/sha_core/w[12] [21]),
	.I1(\top/processor/sha_core/w[13] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_138 )
);
defparam \top/processor/sha_core/n337_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s225  (
	.I0(\top/processor/sha_core/w[14] [21]),
	.I1(\top/processor/sha_core/w[15] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_139 )
);
defparam \top/processor/sha_core/n337_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s226  (
	.I0(\top/processor/sha_core/w[16] [21]),
	.I1(\top/processor/sha_core/w[17] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_140 )
);
defparam \top/processor/sha_core/n337_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s227  (
	.I0(\top/processor/sha_core/w[18] [21]),
	.I1(\top/processor/sha_core/w[19] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_141 )
);
defparam \top/processor/sha_core/n337_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s228  (
	.I0(\top/processor/sha_core/w[20] [21]),
	.I1(\top/processor/sha_core/w[21] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_142 )
);
defparam \top/processor/sha_core/n337_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s229  (
	.I0(\top/processor/sha_core/w[22] [21]),
	.I1(\top/processor/sha_core/w[23] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_143 )
);
defparam \top/processor/sha_core/n337_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s230  (
	.I0(\top/processor/sha_core/w[24] [21]),
	.I1(\top/processor/sha_core/w[25] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_144 )
);
defparam \top/processor/sha_core/n337_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s231  (
	.I0(\top/processor/sha_core/w[26] [21]),
	.I1(\top/processor/sha_core/w[27] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_145 )
);
defparam \top/processor/sha_core/n337_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s232  (
	.I0(\top/processor/sha_core/w[28] [21]),
	.I1(\top/processor/sha_core/w[29] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_146 )
);
defparam \top/processor/sha_core/n337_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s233  (
	.I0(\top/processor/sha_core/w[30] [21]),
	.I1(\top/processor/sha_core/w[31] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_147 )
);
defparam \top/processor/sha_core/n337_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s234  (
	.I0(\top/processor/sha_core/w[32] [21]),
	.I1(\top/processor/sha_core/w[33] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_148 )
);
defparam \top/processor/sha_core/n337_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s235  (
	.I0(\top/processor/sha_core/w[34] [21]),
	.I1(\top/processor/sha_core/w[35] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_149 )
);
defparam \top/processor/sha_core/n337_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s236  (
	.I0(\top/processor/sha_core/w[36] [21]),
	.I1(\top/processor/sha_core/w[37] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_150 )
);
defparam \top/processor/sha_core/n337_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s237  (
	.I0(\top/processor/sha_core/w[38] [21]),
	.I1(\top/processor/sha_core/w[39] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_151 )
);
defparam \top/processor/sha_core/n337_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s238  (
	.I0(\top/processor/sha_core/w[40] [21]),
	.I1(\top/processor/sha_core/w[41] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_152 )
);
defparam \top/processor/sha_core/n337_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s239  (
	.I0(\top/processor/sha_core/w[42] [21]),
	.I1(\top/processor/sha_core/w[43] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_153 )
);
defparam \top/processor/sha_core/n337_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s240  (
	.I0(\top/processor/sha_core/w[44] [21]),
	.I1(\top/processor/sha_core/w[45] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_154 )
);
defparam \top/processor/sha_core/n337_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s241  (
	.I0(\top/processor/sha_core/w[46] [21]),
	.I1(\top/processor/sha_core/w[47] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_155 )
);
defparam \top/processor/sha_core/n337_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s242  (
	.I0(\top/processor/sha_core/w[48] [21]),
	.I1(\top/processor/sha_core/w[49] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_156 )
);
defparam \top/processor/sha_core/n337_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s243  (
	.I0(\top/processor/sha_core/w[50] [21]),
	.I1(\top/processor/sha_core/w[51] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_157 )
);
defparam \top/processor/sha_core/n337_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s244  (
	.I0(\top/processor/sha_core/w[52] [21]),
	.I1(\top/processor/sha_core/w[53] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_158 )
);
defparam \top/processor/sha_core/n337_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s245  (
	.I0(\top/processor/sha_core/w[54] [21]),
	.I1(\top/processor/sha_core/w[55] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_159 )
);
defparam \top/processor/sha_core/n337_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s246  (
	.I0(\top/processor/sha_core/w[56] [21]),
	.I1(\top/processor/sha_core/w[57] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_160 )
);
defparam \top/processor/sha_core/n337_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s247  (
	.I0(\top/processor/sha_core/w[58] [21]),
	.I1(\top/processor/sha_core/w[59] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_161 )
);
defparam \top/processor/sha_core/n337_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s248  (
	.I0(\top/processor/sha_core/w[60] [21]),
	.I1(\top/processor/sha_core/w[61] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_162 )
);
defparam \top/processor/sha_core/n337_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s249  (
	.I0(\top/processor/sha_core/w[62] [21]),
	.I1(\top/processor/sha_core/w[63] [21]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n337_163 )
);
defparam \top/processor/sha_core/n337_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s218  (
	.I0(\top/processor/sha_core/w[0] [20]),
	.I1(\top/processor/sha_core/w[1] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_132 )
);
defparam \top/processor/sha_core/n338_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s219  (
	.I0(\top/processor/sha_core/w[2] [20]),
	.I1(\top/processor/sha_core/w[3] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_133 )
);
defparam \top/processor/sha_core/n338_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s220  (
	.I0(\top/processor/sha_core/w[4] [20]),
	.I1(\top/processor/sha_core/w[5] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_134 )
);
defparam \top/processor/sha_core/n338_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s221  (
	.I0(\top/processor/sha_core/w[6] [20]),
	.I1(\top/processor/sha_core/w[7] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_135 )
);
defparam \top/processor/sha_core/n338_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s222  (
	.I0(\top/processor/sha_core/w[8] [20]),
	.I1(\top/processor/sha_core/w[9] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_136 )
);
defparam \top/processor/sha_core/n338_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s223  (
	.I0(\top/processor/sha_core/w[10] [20]),
	.I1(\top/processor/sha_core/w[11] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_137 )
);
defparam \top/processor/sha_core/n338_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s224  (
	.I0(\top/processor/sha_core/w[12] [20]),
	.I1(\top/processor/sha_core/w[13] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_138 )
);
defparam \top/processor/sha_core/n338_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s225  (
	.I0(\top/processor/sha_core/w[14] [20]),
	.I1(\top/processor/sha_core/w[15] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_139 )
);
defparam \top/processor/sha_core/n338_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s226  (
	.I0(\top/processor/sha_core/w[16] [20]),
	.I1(\top/processor/sha_core/w[17] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_140 )
);
defparam \top/processor/sha_core/n338_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s227  (
	.I0(\top/processor/sha_core/w[18] [20]),
	.I1(\top/processor/sha_core/w[19] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_141 )
);
defparam \top/processor/sha_core/n338_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s228  (
	.I0(\top/processor/sha_core/w[20] [20]),
	.I1(\top/processor/sha_core/w[21] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_142 )
);
defparam \top/processor/sha_core/n338_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s229  (
	.I0(\top/processor/sha_core/w[22] [20]),
	.I1(\top/processor/sha_core/w[23] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_143 )
);
defparam \top/processor/sha_core/n338_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s230  (
	.I0(\top/processor/sha_core/w[24] [20]),
	.I1(\top/processor/sha_core/w[25] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_144 )
);
defparam \top/processor/sha_core/n338_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s231  (
	.I0(\top/processor/sha_core/w[26] [20]),
	.I1(\top/processor/sha_core/w[27] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_145 )
);
defparam \top/processor/sha_core/n338_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s232  (
	.I0(\top/processor/sha_core/w[28] [20]),
	.I1(\top/processor/sha_core/w[29] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_146 )
);
defparam \top/processor/sha_core/n338_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s233  (
	.I0(\top/processor/sha_core/w[30] [20]),
	.I1(\top/processor/sha_core/w[31] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_147 )
);
defparam \top/processor/sha_core/n338_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s234  (
	.I0(\top/processor/sha_core/w[32] [20]),
	.I1(\top/processor/sha_core/w[33] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_148 )
);
defparam \top/processor/sha_core/n338_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s235  (
	.I0(\top/processor/sha_core/w[34] [20]),
	.I1(\top/processor/sha_core/w[35] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_149 )
);
defparam \top/processor/sha_core/n338_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s236  (
	.I0(\top/processor/sha_core/w[36] [20]),
	.I1(\top/processor/sha_core/w[37] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_150 )
);
defparam \top/processor/sha_core/n338_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s237  (
	.I0(\top/processor/sha_core/w[38] [20]),
	.I1(\top/processor/sha_core/w[39] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_151 )
);
defparam \top/processor/sha_core/n338_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s238  (
	.I0(\top/processor/sha_core/w[40] [20]),
	.I1(\top/processor/sha_core/w[41] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_152 )
);
defparam \top/processor/sha_core/n338_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s239  (
	.I0(\top/processor/sha_core/w[42] [20]),
	.I1(\top/processor/sha_core/w[43] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_153 )
);
defparam \top/processor/sha_core/n338_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s240  (
	.I0(\top/processor/sha_core/w[44] [20]),
	.I1(\top/processor/sha_core/w[45] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_154 )
);
defparam \top/processor/sha_core/n338_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s241  (
	.I0(\top/processor/sha_core/w[46] [20]),
	.I1(\top/processor/sha_core/w[47] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_155 )
);
defparam \top/processor/sha_core/n338_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s242  (
	.I0(\top/processor/sha_core/w[48] [20]),
	.I1(\top/processor/sha_core/w[49] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_156 )
);
defparam \top/processor/sha_core/n338_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s243  (
	.I0(\top/processor/sha_core/w[50] [20]),
	.I1(\top/processor/sha_core/w[51] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_157 )
);
defparam \top/processor/sha_core/n338_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s244  (
	.I0(\top/processor/sha_core/w[52] [20]),
	.I1(\top/processor/sha_core/w[53] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_158 )
);
defparam \top/processor/sha_core/n338_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s245  (
	.I0(\top/processor/sha_core/w[54] [20]),
	.I1(\top/processor/sha_core/w[55] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_159 )
);
defparam \top/processor/sha_core/n338_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s246  (
	.I0(\top/processor/sha_core/w[56] [20]),
	.I1(\top/processor/sha_core/w[57] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_160 )
);
defparam \top/processor/sha_core/n338_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s247  (
	.I0(\top/processor/sha_core/w[58] [20]),
	.I1(\top/processor/sha_core/w[59] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_161 )
);
defparam \top/processor/sha_core/n338_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s248  (
	.I0(\top/processor/sha_core/w[60] [20]),
	.I1(\top/processor/sha_core/w[61] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_162 )
);
defparam \top/processor/sha_core/n338_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s249  (
	.I0(\top/processor/sha_core/w[62] [20]),
	.I1(\top/processor/sha_core/w[63] [20]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n338_163 )
);
defparam \top/processor/sha_core/n338_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s218  (
	.I0(\top/processor/sha_core/w[0] [19]),
	.I1(\top/processor/sha_core/w[1] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_132 )
);
defparam \top/processor/sha_core/n339_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s219  (
	.I0(\top/processor/sha_core/w[2] [19]),
	.I1(\top/processor/sha_core/w[3] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_133 )
);
defparam \top/processor/sha_core/n339_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s220  (
	.I0(\top/processor/sha_core/w[4] [19]),
	.I1(\top/processor/sha_core/w[5] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_134 )
);
defparam \top/processor/sha_core/n339_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s221  (
	.I0(\top/processor/sha_core/w[6] [19]),
	.I1(\top/processor/sha_core/w[7] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_135 )
);
defparam \top/processor/sha_core/n339_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s222  (
	.I0(\top/processor/sha_core/w[8] [19]),
	.I1(\top/processor/sha_core/w[9] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_136 )
);
defparam \top/processor/sha_core/n339_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s223  (
	.I0(\top/processor/sha_core/w[10] [19]),
	.I1(\top/processor/sha_core/w[11] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_137 )
);
defparam \top/processor/sha_core/n339_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s224  (
	.I0(\top/processor/sha_core/w[12] [19]),
	.I1(\top/processor/sha_core/w[13] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_138 )
);
defparam \top/processor/sha_core/n339_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s225  (
	.I0(\top/processor/sha_core/w[14] [19]),
	.I1(\top/processor/sha_core/w[15] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_139 )
);
defparam \top/processor/sha_core/n339_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s226  (
	.I0(\top/processor/sha_core/w[16] [19]),
	.I1(\top/processor/sha_core/w[17] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_140 )
);
defparam \top/processor/sha_core/n339_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s227  (
	.I0(\top/processor/sha_core/w[18] [19]),
	.I1(\top/processor/sha_core/w[19] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_141 )
);
defparam \top/processor/sha_core/n339_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s228  (
	.I0(\top/processor/sha_core/w[20] [19]),
	.I1(\top/processor/sha_core/w[21] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_142 )
);
defparam \top/processor/sha_core/n339_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s229  (
	.I0(\top/processor/sha_core/w[22] [19]),
	.I1(\top/processor/sha_core/w[23] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_143 )
);
defparam \top/processor/sha_core/n339_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s230  (
	.I0(\top/processor/sha_core/w[24] [19]),
	.I1(\top/processor/sha_core/w[25] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_144 )
);
defparam \top/processor/sha_core/n339_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s231  (
	.I0(\top/processor/sha_core/w[26] [19]),
	.I1(\top/processor/sha_core/w[27] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_145 )
);
defparam \top/processor/sha_core/n339_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s232  (
	.I0(\top/processor/sha_core/w[28] [19]),
	.I1(\top/processor/sha_core/w[29] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_146 )
);
defparam \top/processor/sha_core/n339_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s233  (
	.I0(\top/processor/sha_core/w[30] [19]),
	.I1(\top/processor/sha_core/w[31] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_147 )
);
defparam \top/processor/sha_core/n339_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s234  (
	.I0(\top/processor/sha_core/w[32] [19]),
	.I1(\top/processor/sha_core/w[33] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_148 )
);
defparam \top/processor/sha_core/n339_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s235  (
	.I0(\top/processor/sha_core/w[34] [19]),
	.I1(\top/processor/sha_core/w[35] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_149 )
);
defparam \top/processor/sha_core/n339_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s236  (
	.I0(\top/processor/sha_core/w[36] [19]),
	.I1(\top/processor/sha_core/w[37] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_150 )
);
defparam \top/processor/sha_core/n339_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s237  (
	.I0(\top/processor/sha_core/w[38] [19]),
	.I1(\top/processor/sha_core/w[39] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_151 )
);
defparam \top/processor/sha_core/n339_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s238  (
	.I0(\top/processor/sha_core/w[40] [19]),
	.I1(\top/processor/sha_core/w[41] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_152 )
);
defparam \top/processor/sha_core/n339_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s239  (
	.I0(\top/processor/sha_core/w[42] [19]),
	.I1(\top/processor/sha_core/w[43] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_153 )
);
defparam \top/processor/sha_core/n339_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s240  (
	.I0(\top/processor/sha_core/w[44] [19]),
	.I1(\top/processor/sha_core/w[45] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_154 )
);
defparam \top/processor/sha_core/n339_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s241  (
	.I0(\top/processor/sha_core/w[46] [19]),
	.I1(\top/processor/sha_core/w[47] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_155 )
);
defparam \top/processor/sha_core/n339_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s242  (
	.I0(\top/processor/sha_core/w[48] [19]),
	.I1(\top/processor/sha_core/w[49] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_156 )
);
defparam \top/processor/sha_core/n339_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s243  (
	.I0(\top/processor/sha_core/w[50] [19]),
	.I1(\top/processor/sha_core/w[51] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_157 )
);
defparam \top/processor/sha_core/n339_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s244  (
	.I0(\top/processor/sha_core/w[52] [19]),
	.I1(\top/processor/sha_core/w[53] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_158 )
);
defparam \top/processor/sha_core/n339_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s245  (
	.I0(\top/processor/sha_core/w[54] [19]),
	.I1(\top/processor/sha_core/w[55] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_159 )
);
defparam \top/processor/sha_core/n339_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s246  (
	.I0(\top/processor/sha_core/w[56] [19]),
	.I1(\top/processor/sha_core/w[57] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_160 )
);
defparam \top/processor/sha_core/n339_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s247  (
	.I0(\top/processor/sha_core/w[58] [19]),
	.I1(\top/processor/sha_core/w[59] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_161 )
);
defparam \top/processor/sha_core/n339_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s248  (
	.I0(\top/processor/sha_core/w[60] [19]),
	.I1(\top/processor/sha_core/w[61] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_162 )
);
defparam \top/processor/sha_core/n339_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s249  (
	.I0(\top/processor/sha_core/w[62] [19]),
	.I1(\top/processor/sha_core/w[63] [19]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n339_163 )
);
defparam \top/processor/sha_core/n339_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s218  (
	.I0(\top/processor/sha_core/w[0] [18]),
	.I1(\top/processor/sha_core/w[1] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_132 )
);
defparam \top/processor/sha_core/n340_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s219  (
	.I0(\top/processor/sha_core/w[2] [18]),
	.I1(\top/processor/sha_core/w[3] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_133 )
);
defparam \top/processor/sha_core/n340_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s220  (
	.I0(\top/processor/sha_core/w[4] [18]),
	.I1(\top/processor/sha_core/w[5] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_134 )
);
defparam \top/processor/sha_core/n340_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s221  (
	.I0(\top/processor/sha_core/w[6] [18]),
	.I1(\top/processor/sha_core/w[7] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_135 )
);
defparam \top/processor/sha_core/n340_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s222  (
	.I0(\top/processor/sha_core/w[8] [18]),
	.I1(\top/processor/sha_core/w[9] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_136 )
);
defparam \top/processor/sha_core/n340_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s223  (
	.I0(\top/processor/sha_core/w[10] [18]),
	.I1(\top/processor/sha_core/w[11] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_137 )
);
defparam \top/processor/sha_core/n340_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s224  (
	.I0(\top/processor/sha_core/w[12] [18]),
	.I1(\top/processor/sha_core/w[13] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_138 )
);
defparam \top/processor/sha_core/n340_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s225  (
	.I0(\top/processor/sha_core/w[14] [18]),
	.I1(\top/processor/sha_core/w[15] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_139 )
);
defparam \top/processor/sha_core/n340_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s226  (
	.I0(\top/processor/sha_core/w[16] [18]),
	.I1(\top/processor/sha_core/w[17] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_140 )
);
defparam \top/processor/sha_core/n340_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s227  (
	.I0(\top/processor/sha_core/w[18] [18]),
	.I1(\top/processor/sha_core/w[19] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_141 )
);
defparam \top/processor/sha_core/n340_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s228  (
	.I0(\top/processor/sha_core/w[20] [18]),
	.I1(\top/processor/sha_core/w[21] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_142 )
);
defparam \top/processor/sha_core/n340_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s229  (
	.I0(\top/processor/sha_core/w[22] [18]),
	.I1(\top/processor/sha_core/w[23] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_143 )
);
defparam \top/processor/sha_core/n340_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s230  (
	.I0(\top/processor/sha_core/w[24] [18]),
	.I1(\top/processor/sha_core/w[25] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_144 )
);
defparam \top/processor/sha_core/n340_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s231  (
	.I0(\top/processor/sha_core/w[26] [18]),
	.I1(\top/processor/sha_core/w[27] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_145 )
);
defparam \top/processor/sha_core/n340_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s232  (
	.I0(\top/processor/sha_core/w[28] [18]),
	.I1(\top/processor/sha_core/w[29] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_146 )
);
defparam \top/processor/sha_core/n340_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s233  (
	.I0(\top/processor/sha_core/w[30] [18]),
	.I1(\top/processor/sha_core/w[31] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_147 )
);
defparam \top/processor/sha_core/n340_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s234  (
	.I0(\top/processor/sha_core/w[32] [18]),
	.I1(\top/processor/sha_core/w[33] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_148 )
);
defparam \top/processor/sha_core/n340_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s235  (
	.I0(\top/processor/sha_core/w[34] [18]),
	.I1(\top/processor/sha_core/w[35] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_149 )
);
defparam \top/processor/sha_core/n340_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s236  (
	.I0(\top/processor/sha_core/w[36] [18]),
	.I1(\top/processor/sha_core/w[37] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_150 )
);
defparam \top/processor/sha_core/n340_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s237  (
	.I0(\top/processor/sha_core/w[38] [18]),
	.I1(\top/processor/sha_core/w[39] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_151 )
);
defparam \top/processor/sha_core/n340_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s238  (
	.I0(\top/processor/sha_core/w[40] [18]),
	.I1(\top/processor/sha_core/w[41] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_152 )
);
defparam \top/processor/sha_core/n340_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s239  (
	.I0(\top/processor/sha_core/w[42] [18]),
	.I1(\top/processor/sha_core/w[43] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_153 )
);
defparam \top/processor/sha_core/n340_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s240  (
	.I0(\top/processor/sha_core/w[44] [18]),
	.I1(\top/processor/sha_core/w[45] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_154 )
);
defparam \top/processor/sha_core/n340_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s241  (
	.I0(\top/processor/sha_core/w[46] [18]),
	.I1(\top/processor/sha_core/w[47] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_155 )
);
defparam \top/processor/sha_core/n340_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s242  (
	.I0(\top/processor/sha_core/w[48] [18]),
	.I1(\top/processor/sha_core/w[49] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_156 )
);
defparam \top/processor/sha_core/n340_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s243  (
	.I0(\top/processor/sha_core/w[50] [18]),
	.I1(\top/processor/sha_core/w[51] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_157 )
);
defparam \top/processor/sha_core/n340_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s244  (
	.I0(\top/processor/sha_core/w[52] [18]),
	.I1(\top/processor/sha_core/w[53] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_158 )
);
defparam \top/processor/sha_core/n340_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s245  (
	.I0(\top/processor/sha_core/w[54] [18]),
	.I1(\top/processor/sha_core/w[55] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_159 )
);
defparam \top/processor/sha_core/n340_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s246  (
	.I0(\top/processor/sha_core/w[56] [18]),
	.I1(\top/processor/sha_core/w[57] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_160 )
);
defparam \top/processor/sha_core/n340_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s247  (
	.I0(\top/processor/sha_core/w[58] [18]),
	.I1(\top/processor/sha_core/w[59] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_161 )
);
defparam \top/processor/sha_core/n340_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s248  (
	.I0(\top/processor/sha_core/w[60] [18]),
	.I1(\top/processor/sha_core/w[61] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_162 )
);
defparam \top/processor/sha_core/n340_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s249  (
	.I0(\top/processor/sha_core/w[62] [18]),
	.I1(\top/processor/sha_core/w[63] [18]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n340_163 )
);
defparam \top/processor/sha_core/n340_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s218  (
	.I0(\top/processor/sha_core/w[0] [17]),
	.I1(\top/processor/sha_core/w[1] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_132 )
);
defparam \top/processor/sha_core/n341_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s219  (
	.I0(\top/processor/sha_core/w[2] [17]),
	.I1(\top/processor/sha_core/w[3] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_133 )
);
defparam \top/processor/sha_core/n341_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s220  (
	.I0(\top/processor/sha_core/w[4] [17]),
	.I1(\top/processor/sha_core/w[5] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_134 )
);
defparam \top/processor/sha_core/n341_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s221  (
	.I0(\top/processor/sha_core/w[6] [17]),
	.I1(\top/processor/sha_core/w[7] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_135 )
);
defparam \top/processor/sha_core/n341_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s222  (
	.I0(\top/processor/sha_core/w[8] [17]),
	.I1(\top/processor/sha_core/w[9] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_136 )
);
defparam \top/processor/sha_core/n341_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s223  (
	.I0(\top/processor/sha_core/w[10] [17]),
	.I1(\top/processor/sha_core/w[11] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_137 )
);
defparam \top/processor/sha_core/n341_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s224  (
	.I0(\top/processor/sha_core/w[12] [17]),
	.I1(\top/processor/sha_core/w[13] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_138 )
);
defparam \top/processor/sha_core/n341_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s225  (
	.I0(\top/processor/sha_core/w[14] [17]),
	.I1(\top/processor/sha_core/w[15] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_139 )
);
defparam \top/processor/sha_core/n341_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s226  (
	.I0(\top/processor/sha_core/w[16] [17]),
	.I1(\top/processor/sha_core/w[17] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_140 )
);
defparam \top/processor/sha_core/n341_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s227  (
	.I0(\top/processor/sha_core/w[18] [17]),
	.I1(\top/processor/sha_core/w[19] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_141 )
);
defparam \top/processor/sha_core/n341_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s228  (
	.I0(\top/processor/sha_core/w[20] [17]),
	.I1(\top/processor/sha_core/w[21] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_142 )
);
defparam \top/processor/sha_core/n341_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s229  (
	.I0(\top/processor/sha_core/w[22] [17]),
	.I1(\top/processor/sha_core/w[23] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_143 )
);
defparam \top/processor/sha_core/n341_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s230  (
	.I0(\top/processor/sha_core/w[24] [17]),
	.I1(\top/processor/sha_core/w[25] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_144 )
);
defparam \top/processor/sha_core/n341_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s231  (
	.I0(\top/processor/sha_core/w[26] [17]),
	.I1(\top/processor/sha_core/w[27] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_145 )
);
defparam \top/processor/sha_core/n341_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s232  (
	.I0(\top/processor/sha_core/w[28] [17]),
	.I1(\top/processor/sha_core/w[29] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_146 )
);
defparam \top/processor/sha_core/n341_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s233  (
	.I0(\top/processor/sha_core/w[30] [17]),
	.I1(\top/processor/sha_core/w[31] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_147 )
);
defparam \top/processor/sha_core/n341_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s234  (
	.I0(\top/processor/sha_core/w[32] [17]),
	.I1(\top/processor/sha_core/w[33] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_148 )
);
defparam \top/processor/sha_core/n341_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s235  (
	.I0(\top/processor/sha_core/w[34] [17]),
	.I1(\top/processor/sha_core/w[35] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_149 )
);
defparam \top/processor/sha_core/n341_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s236  (
	.I0(\top/processor/sha_core/w[36] [17]),
	.I1(\top/processor/sha_core/w[37] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_150 )
);
defparam \top/processor/sha_core/n341_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s237  (
	.I0(\top/processor/sha_core/w[38] [17]),
	.I1(\top/processor/sha_core/w[39] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_151 )
);
defparam \top/processor/sha_core/n341_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s238  (
	.I0(\top/processor/sha_core/w[40] [17]),
	.I1(\top/processor/sha_core/w[41] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_152 )
);
defparam \top/processor/sha_core/n341_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s239  (
	.I0(\top/processor/sha_core/w[42] [17]),
	.I1(\top/processor/sha_core/w[43] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_153 )
);
defparam \top/processor/sha_core/n341_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s240  (
	.I0(\top/processor/sha_core/w[44] [17]),
	.I1(\top/processor/sha_core/w[45] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_154 )
);
defparam \top/processor/sha_core/n341_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s241  (
	.I0(\top/processor/sha_core/w[46] [17]),
	.I1(\top/processor/sha_core/w[47] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_155 )
);
defparam \top/processor/sha_core/n341_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s242  (
	.I0(\top/processor/sha_core/w[48] [17]),
	.I1(\top/processor/sha_core/w[49] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_156 )
);
defparam \top/processor/sha_core/n341_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s243  (
	.I0(\top/processor/sha_core/w[50] [17]),
	.I1(\top/processor/sha_core/w[51] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_157 )
);
defparam \top/processor/sha_core/n341_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s244  (
	.I0(\top/processor/sha_core/w[52] [17]),
	.I1(\top/processor/sha_core/w[53] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_158 )
);
defparam \top/processor/sha_core/n341_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s245  (
	.I0(\top/processor/sha_core/w[54] [17]),
	.I1(\top/processor/sha_core/w[55] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_159 )
);
defparam \top/processor/sha_core/n341_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s246  (
	.I0(\top/processor/sha_core/w[56] [17]),
	.I1(\top/processor/sha_core/w[57] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_160 )
);
defparam \top/processor/sha_core/n341_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s247  (
	.I0(\top/processor/sha_core/w[58] [17]),
	.I1(\top/processor/sha_core/w[59] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_161 )
);
defparam \top/processor/sha_core/n341_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s248  (
	.I0(\top/processor/sha_core/w[60] [17]),
	.I1(\top/processor/sha_core/w[61] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_162 )
);
defparam \top/processor/sha_core/n341_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s249  (
	.I0(\top/processor/sha_core/w[62] [17]),
	.I1(\top/processor/sha_core/w[63] [17]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n341_163 )
);
defparam \top/processor/sha_core/n341_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s218  (
	.I0(\top/processor/sha_core/w[0] [16]),
	.I1(\top/processor/sha_core/w[1] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_132 )
);
defparam \top/processor/sha_core/n342_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s219  (
	.I0(\top/processor/sha_core/w[2] [16]),
	.I1(\top/processor/sha_core/w[3] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_133 )
);
defparam \top/processor/sha_core/n342_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s220  (
	.I0(\top/processor/sha_core/w[4] [16]),
	.I1(\top/processor/sha_core/w[5] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_134 )
);
defparam \top/processor/sha_core/n342_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s221  (
	.I0(\top/processor/sha_core/w[6] [16]),
	.I1(\top/processor/sha_core/w[7] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_135 )
);
defparam \top/processor/sha_core/n342_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s222  (
	.I0(\top/processor/sha_core/w[8] [16]),
	.I1(\top/processor/sha_core/w[9] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_136 )
);
defparam \top/processor/sha_core/n342_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s223  (
	.I0(\top/processor/sha_core/w[10] [16]),
	.I1(\top/processor/sha_core/w[11] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_137 )
);
defparam \top/processor/sha_core/n342_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s224  (
	.I0(\top/processor/sha_core/w[12] [16]),
	.I1(\top/processor/sha_core/w[13] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_138 )
);
defparam \top/processor/sha_core/n342_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s225  (
	.I0(\top/processor/sha_core/w[14] [16]),
	.I1(\top/processor/sha_core/w[15] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_139 )
);
defparam \top/processor/sha_core/n342_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s226  (
	.I0(\top/processor/sha_core/w[16] [16]),
	.I1(\top/processor/sha_core/w[17] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_140 )
);
defparam \top/processor/sha_core/n342_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s227  (
	.I0(\top/processor/sha_core/w[18] [16]),
	.I1(\top/processor/sha_core/w[19] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_141 )
);
defparam \top/processor/sha_core/n342_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s228  (
	.I0(\top/processor/sha_core/w[20] [16]),
	.I1(\top/processor/sha_core/w[21] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_142 )
);
defparam \top/processor/sha_core/n342_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s229  (
	.I0(\top/processor/sha_core/w[22] [16]),
	.I1(\top/processor/sha_core/w[23] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_143 )
);
defparam \top/processor/sha_core/n342_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s230  (
	.I0(\top/processor/sha_core/w[24] [16]),
	.I1(\top/processor/sha_core/w[25] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_144 )
);
defparam \top/processor/sha_core/n342_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s231  (
	.I0(\top/processor/sha_core/w[26] [16]),
	.I1(\top/processor/sha_core/w[27] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_145 )
);
defparam \top/processor/sha_core/n342_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s232  (
	.I0(\top/processor/sha_core/w[28] [16]),
	.I1(\top/processor/sha_core/w[29] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_146 )
);
defparam \top/processor/sha_core/n342_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s233  (
	.I0(\top/processor/sha_core/w[30] [16]),
	.I1(\top/processor/sha_core/w[31] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_147 )
);
defparam \top/processor/sha_core/n342_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s234  (
	.I0(\top/processor/sha_core/w[32] [16]),
	.I1(\top/processor/sha_core/w[33] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_148 )
);
defparam \top/processor/sha_core/n342_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s235  (
	.I0(\top/processor/sha_core/w[34] [16]),
	.I1(\top/processor/sha_core/w[35] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_149 )
);
defparam \top/processor/sha_core/n342_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s236  (
	.I0(\top/processor/sha_core/w[36] [16]),
	.I1(\top/processor/sha_core/w[37] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_150 )
);
defparam \top/processor/sha_core/n342_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s237  (
	.I0(\top/processor/sha_core/w[38] [16]),
	.I1(\top/processor/sha_core/w[39] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_151 )
);
defparam \top/processor/sha_core/n342_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s238  (
	.I0(\top/processor/sha_core/w[40] [16]),
	.I1(\top/processor/sha_core/w[41] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_152 )
);
defparam \top/processor/sha_core/n342_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s239  (
	.I0(\top/processor/sha_core/w[42] [16]),
	.I1(\top/processor/sha_core/w[43] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_153 )
);
defparam \top/processor/sha_core/n342_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s240  (
	.I0(\top/processor/sha_core/w[44] [16]),
	.I1(\top/processor/sha_core/w[45] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_154 )
);
defparam \top/processor/sha_core/n342_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s241  (
	.I0(\top/processor/sha_core/w[46] [16]),
	.I1(\top/processor/sha_core/w[47] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_155 )
);
defparam \top/processor/sha_core/n342_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s242  (
	.I0(\top/processor/sha_core/w[48] [16]),
	.I1(\top/processor/sha_core/w[49] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_156 )
);
defparam \top/processor/sha_core/n342_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s243  (
	.I0(\top/processor/sha_core/w[50] [16]),
	.I1(\top/processor/sha_core/w[51] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_157 )
);
defparam \top/processor/sha_core/n342_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s244  (
	.I0(\top/processor/sha_core/w[52] [16]),
	.I1(\top/processor/sha_core/w[53] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_158 )
);
defparam \top/processor/sha_core/n342_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s245  (
	.I0(\top/processor/sha_core/w[54] [16]),
	.I1(\top/processor/sha_core/w[55] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_159 )
);
defparam \top/processor/sha_core/n342_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s246  (
	.I0(\top/processor/sha_core/w[56] [16]),
	.I1(\top/processor/sha_core/w[57] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_160 )
);
defparam \top/processor/sha_core/n342_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s247  (
	.I0(\top/processor/sha_core/w[58] [16]),
	.I1(\top/processor/sha_core/w[59] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_161 )
);
defparam \top/processor/sha_core/n342_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s248  (
	.I0(\top/processor/sha_core/w[60] [16]),
	.I1(\top/processor/sha_core/w[61] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_162 )
);
defparam \top/processor/sha_core/n342_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s249  (
	.I0(\top/processor/sha_core/w[62] [16]),
	.I1(\top/processor/sha_core/w[63] [16]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n342_163 )
);
defparam \top/processor/sha_core/n342_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s218  (
	.I0(\top/processor/sha_core/w[0] [15]),
	.I1(\top/processor/sha_core/w[1] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_132 )
);
defparam \top/processor/sha_core/n343_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s219  (
	.I0(\top/processor/sha_core/w[2] [15]),
	.I1(\top/processor/sha_core/w[3] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_133 )
);
defparam \top/processor/sha_core/n343_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s220  (
	.I0(\top/processor/sha_core/w[4] [15]),
	.I1(\top/processor/sha_core/w[5] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_134 )
);
defparam \top/processor/sha_core/n343_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s221  (
	.I0(\top/processor/sha_core/w[6] [15]),
	.I1(\top/processor/sha_core/w[7] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_135 )
);
defparam \top/processor/sha_core/n343_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s222  (
	.I0(\top/processor/sha_core/w[8] [15]),
	.I1(\top/processor/sha_core/w[9] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_136 )
);
defparam \top/processor/sha_core/n343_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s223  (
	.I0(\top/processor/sha_core/w[10] [15]),
	.I1(\top/processor/sha_core/w[11] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_137 )
);
defparam \top/processor/sha_core/n343_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s224  (
	.I0(\top/processor/sha_core/w[12] [15]),
	.I1(\top/processor/sha_core/w[13] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_138 )
);
defparam \top/processor/sha_core/n343_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s225  (
	.I0(\top/processor/sha_core/w[14] [15]),
	.I1(\top/processor/sha_core/w[15] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_139 )
);
defparam \top/processor/sha_core/n343_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s226  (
	.I0(\top/processor/sha_core/w[16] [15]),
	.I1(\top/processor/sha_core/w[17] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_140 )
);
defparam \top/processor/sha_core/n343_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s227  (
	.I0(\top/processor/sha_core/w[18] [15]),
	.I1(\top/processor/sha_core/w[19] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_141 )
);
defparam \top/processor/sha_core/n343_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s228  (
	.I0(\top/processor/sha_core/w[20] [15]),
	.I1(\top/processor/sha_core/w[21] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_142 )
);
defparam \top/processor/sha_core/n343_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s229  (
	.I0(\top/processor/sha_core/w[22] [15]),
	.I1(\top/processor/sha_core/w[23] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_143 )
);
defparam \top/processor/sha_core/n343_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s230  (
	.I0(\top/processor/sha_core/w[24] [15]),
	.I1(\top/processor/sha_core/w[25] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_144 )
);
defparam \top/processor/sha_core/n343_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s231  (
	.I0(\top/processor/sha_core/w[26] [15]),
	.I1(\top/processor/sha_core/w[27] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_145 )
);
defparam \top/processor/sha_core/n343_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s232  (
	.I0(\top/processor/sha_core/w[28] [15]),
	.I1(\top/processor/sha_core/w[29] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_146 )
);
defparam \top/processor/sha_core/n343_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s233  (
	.I0(\top/processor/sha_core/w[30] [15]),
	.I1(\top/processor/sha_core/w[31] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_147 )
);
defparam \top/processor/sha_core/n343_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s234  (
	.I0(\top/processor/sha_core/w[32] [15]),
	.I1(\top/processor/sha_core/w[33] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_148 )
);
defparam \top/processor/sha_core/n343_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s235  (
	.I0(\top/processor/sha_core/w[34] [15]),
	.I1(\top/processor/sha_core/w[35] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_149 )
);
defparam \top/processor/sha_core/n343_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s236  (
	.I0(\top/processor/sha_core/w[36] [15]),
	.I1(\top/processor/sha_core/w[37] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_150 )
);
defparam \top/processor/sha_core/n343_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s237  (
	.I0(\top/processor/sha_core/w[38] [15]),
	.I1(\top/processor/sha_core/w[39] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_151 )
);
defparam \top/processor/sha_core/n343_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s238  (
	.I0(\top/processor/sha_core/w[40] [15]),
	.I1(\top/processor/sha_core/w[41] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_152 )
);
defparam \top/processor/sha_core/n343_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s239  (
	.I0(\top/processor/sha_core/w[42] [15]),
	.I1(\top/processor/sha_core/w[43] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_153 )
);
defparam \top/processor/sha_core/n343_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s240  (
	.I0(\top/processor/sha_core/w[44] [15]),
	.I1(\top/processor/sha_core/w[45] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_154 )
);
defparam \top/processor/sha_core/n343_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s241  (
	.I0(\top/processor/sha_core/w[46] [15]),
	.I1(\top/processor/sha_core/w[47] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_155 )
);
defparam \top/processor/sha_core/n343_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s242  (
	.I0(\top/processor/sha_core/w[48] [15]),
	.I1(\top/processor/sha_core/w[49] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_156 )
);
defparam \top/processor/sha_core/n343_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s243  (
	.I0(\top/processor/sha_core/w[50] [15]),
	.I1(\top/processor/sha_core/w[51] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_157 )
);
defparam \top/processor/sha_core/n343_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s244  (
	.I0(\top/processor/sha_core/w[52] [15]),
	.I1(\top/processor/sha_core/w[53] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_158 )
);
defparam \top/processor/sha_core/n343_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s245  (
	.I0(\top/processor/sha_core/w[54] [15]),
	.I1(\top/processor/sha_core/w[55] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_159 )
);
defparam \top/processor/sha_core/n343_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s246  (
	.I0(\top/processor/sha_core/w[56] [15]),
	.I1(\top/processor/sha_core/w[57] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_160 )
);
defparam \top/processor/sha_core/n343_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s247  (
	.I0(\top/processor/sha_core/w[58] [15]),
	.I1(\top/processor/sha_core/w[59] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_161 )
);
defparam \top/processor/sha_core/n343_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s248  (
	.I0(\top/processor/sha_core/w[60] [15]),
	.I1(\top/processor/sha_core/w[61] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_162 )
);
defparam \top/processor/sha_core/n343_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s249  (
	.I0(\top/processor/sha_core/w[62] [15]),
	.I1(\top/processor/sha_core/w[63] [15]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n343_163 )
);
defparam \top/processor/sha_core/n343_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s218  (
	.I0(\top/processor/sha_core/w[0] [14]),
	.I1(\top/processor/sha_core/w[1] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_132 )
);
defparam \top/processor/sha_core/n344_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s219  (
	.I0(\top/processor/sha_core/w[2] [14]),
	.I1(\top/processor/sha_core/w[3] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_133 )
);
defparam \top/processor/sha_core/n344_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s220  (
	.I0(\top/processor/sha_core/w[4] [14]),
	.I1(\top/processor/sha_core/w[5] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_134 )
);
defparam \top/processor/sha_core/n344_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s221  (
	.I0(\top/processor/sha_core/w[6] [14]),
	.I1(\top/processor/sha_core/w[7] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_135 )
);
defparam \top/processor/sha_core/n344_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s222  (
	.I0(\top/processor/sha_core/w[8] [14]),
	.I1(\top/processor/sha_core/w[9] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_136 )
);
defparam \top/processor/sha_core/n344_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s223  (
	.I0(\top/processor/sha_core/w[10] [14]),
	.I1(\top/processor/sha_core/w[11] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_137 )
);
defparam \top/processor/sha_core/n344_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s224  (
	.I0(\top/processor/sha_core/w[12] [14]),
	.I1(\top/processor/sha_core/w[13] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_138 )
);
defparam \top/processor/sha_core/n344_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s225  (
	.I0(\top/processor/sha_core/w[14] [14]),
	.I1(\top/processor/sha_core/w[15] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_139 )
);
defparam \top/processor/sha_core/n344_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s226  (
	.I0(\top/processor/sha_core/w[16] [14]),
	.I1(\top/processor/sha_core/w[17] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_140 )
);
defparam \top/processor/sha_core/n344_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s227  (
	.I0(\top/processor/sha_core/w[18] [14]),
	.I1(\top/processor/sha_core/w[19] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_141 )
);
defparam \top/processor/sha_core/n344_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s228  (
	.I0(\top/processor/sha_core/w[20] [14]),
	.I1(\top/processor/sha_core/w[21] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_142 )
);
defparam \top/processor/sha_core/n344_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s229  (
	.I0(\top/processor/sha_core/w[22] [14]),
	.I1(\top/processor/sha_core/w[23] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_143 )
);
defparam \top/processor/sha_core/n344_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s230  (
	.I0(\top/processor/sha_core/w[24] [14]),
	.I1(\top/processor/sha_core/w[25] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_144 )
);
defparam \top/processor/sha_core/n344_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s231  (
	.I0(\top/processor/sha_core/w[26] [14]),
	.I1(\top/processor/sha_core/w[27] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_145 )
);
defparam \top/processor/sha_core/n344_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s232  (
	.I0(\top/processor/sha_core/w[28] [14]),
	.I1(\top/processor/sha_core/w[29] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_146 )
);
defparam \top/processor/sha_core/n344_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s233  (
	.I0(\top/processor/sha_core/w[30] [14]),
	.I1(\top/processor/sha_core/w[31] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_147 )
);
defparam \top/processor/sha_core/n344_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s234  (
	.I0(\top/processor/sha_core/w[32] [14]),
	.I1(\top/processor/sha_core/w[33] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_148 )
);
defparam \top/processor/sha_core/n344_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s235  (
	.I0(\top/processor/sha_core/w[34] [14]),
	.I1(\top/processor/sha_core/w[35] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_149 )
);
defparam \top/processor/sha_core/n344_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s236  (
	.I0(\top/processor/sha_core/w[36] [14]),
	.I1(\top/processor/sha_core/w[37] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_150 )
);
defparam \top/processor/sha_core/n344_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s237  (
	.I0(\top/processor/sha_core/w[38] [14]),
	.I1(\top/processor/sha_core/w[39] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_151 )
);
defparam \top/processor/sha_core/n344_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s238  (
	.I0(\top/processor/sha_core/w[40] [14]),
	.I1(\top/processor/sha_core/w[41] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_152 )
);
defparam \top/processor/sha_core/n344_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s239  (
	.I0(\top/processor/sha_core/w[42] [14]),
	.I1(\top/processor/sha_core/w[43] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_153 )
);
defparam \top/processor/sha_core/n344_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s240  (
	.I0(\top/processor/sha_core/w[44] [14]),
	.I1(\top/processor/sha_core/w[45] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_154 )
);
defparam \top/processor/sha_core/n344_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s241  (
	.I0(\top/processor/sha_core/w[46] [14]),
	.I1(\top/processor/sha_core/w[47] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_155 )
);
defparam \top/processor/sha_core/n344_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s242  (
	.I0(\top/processor/sha_core/w[48] [14]),
	.I1(\top/processor/sha_core/w[49] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_156 )
);
defparam \top/processor/sha_core/n344_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s243  (
	.I0(\top/processor/sha_core/w[50] [14]),
	.I1(\top/processor/sha_core/w[51] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_157 )
);
defparam \top/processor/sha_core/n344_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s244  (
	.I0(\top/processor/sha_core/w[52] [14]),
	.I1(\top/processor/sha_core/w[53] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_158 )
);
defparam \top/processor/sha_core/n344_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s245  (
	.I0(\top/processor/sha_core/w[54] [14]),
	.I1(\top/processor/sha_core/w[55] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_159 )
);
defparam \top/processor/sha_core/n344_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s246  (
	.I0(\top/processor/sha_core/w[56] [14]),
	.I1(\top/processor/sha_core/w[57] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_160 )
);
defparam \top/processor/sha_core/n344_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s247  (
	.I0(\top/processor/sha_core/w[58] [14]),
	.I1(\top/processor/sha_core/w[59] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_161 )
);
defparam \top/processor/sha_core/n344_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s248  (
	.I0(\top/processor/sha_core/w[60] [14]),
	.I1(\top/processor/sha_core/w[61] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_162 )
);
defparam \top/processor/sha_core/n344_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s249  (
	.I0(\top/processor/sha_core/w[62] [14]),
	.I1(\top/processor/sha_core/w[63] [14]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n344_163 )
);
defparam \top/processor/sha_core/n344_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s218  (
	.I0(\top/processor/sha_core/w[0] [13]),
	.I1(\top/processor/sha_core/w[1] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_132 )
);
defparam \top/processor/sha_core/n345_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s219  (
	.I0(\top/processor/sha_core/w[2] [13]),
	.I1(\top/processor/sha_core/w[3] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_133 )
);
defparam \top/processor/sha_core/n345_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s220  (
	.I0(\top/processor/sha_core/w[4] [13]),
	.I1(\top/processor/sha_core/w[5] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_134 )
);
defparam \top/processor/sha_core/n345_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s221  (
	.I0(\top/processor/sha_core/w[6] [13]),
	.I1(\top/processor/sha_core/w[7] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_135 )
);
defparam \top/processor/sha_core/n345_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s222  (
	.I0(\top/processor/sha_core/w[8] [13]),
	.I1(\top/processor/sha_core/w[9] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_136 )
);
defparam \top/processor/sha_core/n345_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s223  (
	.I0(\top/processor/sha_core/w[10] [13]),
	.I1(\top/processor/sha_core/w[11] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_137 )
);
defparam \top/processor/sha_core/n345_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s224  (
	.I0(\top/processor/sha_core/w[12] [13]),
	.I1(\top/processor/sha_core/w[13] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_138 )
);
defparam \top/processor/sha_core/n345_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s225  (
	.I0(\top/processor/sha_core/w[14] [13]),
	.I1(\top/processor/sha_core/w[15] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_139 )
);
defparam \top/processor/sha_core/n345_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s226  (
	.I0(\top/processor/sha_core/w[16] [13]),
	.I1(\top/processor/sha_core/w[17] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_140 )
);
defparam \top/processor/sha_core/n345_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s227  (
	.I0(\top/processor/sha_core/w[18] [13]),
	.I1(\top/processor/sha_core/w[19] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_141 )
);
defparam \top/processor/sha_core/n345_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s228  (
	.I0(\top/processor/sha_core/w[20] [13]),
	.I1(\top/processor/sha_core/w[21] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_142 )
);
defparam \top/processor/sha_core/n345_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s229  (
	.I0(\top/processor/sha_core/w[22] [13]),
	.I1(\top/processor/sha_core/w[23] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_143 )
);
defparam \top/processor/sha_core/n345_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s230  (
	.I0(\top/processor/sha_core/w[24] [13]),
	.I1(\top/processor/sha_core/w[25] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_144 )
);
defparam \top/processor/sha_core/n345_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s231  (
	.I0(\top/processor/sha_core/w[26] [13]),
	.I1(\top/processor/sha_core/w[27] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_145 )
);
defparam \top/processor/sha_core/n345_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s232  (
	.I0(\top/processor/sha_core/w[28] [13]),
	.I1(\top/processor/sha_core/w[29] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_146 )
);
defparam \top/processor/sha_core/n345_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s233  (
	.I0(\top/processor/sha_core/w[30] [13]),
	.I1(\top/processor/sha_core/w[31] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_147 )
);
defparam \top/processor/sha_core/n345_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s234  (
	.I0(\top/processor/sha_core/w[32] [13]),
	.I1(\top/processor/sha_core/w[33] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_148 )
);
defparam \top/processor/sha_core/n345_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s235  (
	.I0(\top/processor/sha_core/w[34] [13]),
	.I1(\top/processor/sha_core/w[35] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_149 )
);
defparam \top/processor/sha_core/n345_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s236  (
	.I0(\top/processor/sha_core/w[36] [13]),
	.I1(\top/processor/sha_core/w[37] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_150 )
);
defparam \top/processor/sha_core/n345_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s237  (
	.I0(\top/processor/sha_core/w[38] [13]),
	.I1(\top/processor/sha_core/w[39] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_151 )
);
defparam \top/processor/sha_core/n345_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s238  (
	.I0(\top/processor/sha_core/w[40] [13]),
	.I1(\top/processor/sha_core/w[41] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_152 )
);
defparam \top/processor/sha_core/n345_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s239  (
	.I0(\top/processor/sha_core/w[42] [13]),
	.I1(\top/processor/sha_core/w[43] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_153 )
);
defparam \top/processor/sha_core/n345_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s240  (
	.I0(\top/processor/sha_core/w[44] [13]),
	.I1(\top/processor/sha_core/w[45] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_154 )
);
defparam \top/processor/sha_core/n345_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s241  (
	.I0(\top/processor/sha_core/w[46] [13]),
	.I1(\top/processor/sha_core/w[47] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_155 )
);
defparam \top/processor/sha_core/n345_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s242  (
	.I0(\top/processor/sha_core/w[48] [13]),
	.I1(\top/processor/sha_core/w[49] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_156 )
);
defparam \top/processor/sha_core/n345_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s243  (
	.I0(\top/processor/sha_core/w[50] [13]),
	.I1(\top/processor/sha_core/w[51] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_157 )
);
defparam \top/processor/sha_core/n345_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s244  (
	.I0(\top/processor/sha_core/w[52] [13]),
	.I1(\top/processor/sha_core/w[53] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_158 )
);
defparam \top/processor/sha_core/n345_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s245  (
	.I0(\top/processor/sha_core/w[54] [13]),
	.I1(\top/processor/sha_core/w[55] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_159 )
);
defparam \top/processor/sha_core/n345_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s246  (
	.I0(\top/processor/sha_core/w[56] [13]),
	.I1(\top/processor/sha_core/w[57] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_160 )
);
defparam \top/processor/sha_core/n345_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s247  (
	.I0(\top/processor/sha_core/w[58] [13]),
	.I1(\top/processor/sha_core/w[59] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_161 )
);
defparam \top/processor/sha_core/n345_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s248  (
	.I0(\top/processor/sha_core/w[60] [13]),
	.I1(\top/processor/sha_core/w[61] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_162 )
);
defparam \top/processor/sha_core/n345_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s249  (
	.I0(\top/processor/sha_core/w[62] [13]),
	.I1(\top/processor/sha_core/w[63] [13]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n345_163 )
);
defparam \top/processor/sha_core/n345_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s218  (
	.I0(\top/processor/sha_core/w[0] [12]),
	.I1(\top/processor/sha_core/w[1] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_132 )
);
defparam \top/processor/sha_core/n346_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s219  (
	.I0(\top/processor/sha_core/w[2] [12]),
	.I1(\top/processor/sha_core/w[3] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_133 )
);
defparam \top/processor/sha_core/n346_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s220  (
	.I0(\top/processor/sha_core/w[4] [12]),
	.I1(\top/processor/sha_core/w[5] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_134 )
);
defparam \top/processor/sha_core/n346_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s221  (
	.I0(\top/processor/sha_core/w[6] [12]),
	.I1(\top/processor/sha_core/w[7] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_135 )
);
defparam \top/processor/sha_core/n346_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s222  (
	.I0(\top/processor/sha_core/w[8] [12]),
	.I1(\top/processor/sha_core/w[9] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_136 )
);
defparam \top/processor/sha_core/n346_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s223  (
	.I0(\top/processor/sha_core/w[10] [12]),
	.I1(\top/processor/sha_core/w[11] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_137 )
);
defparam \top/processor/sha_core/n346_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s224  (
	.I0(\top/processor/sha_core/w[12] [12]),
	.I1(\top/processor/sha_core/w[13] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_138 )
);
defparam \top/processor/sha_core/n346_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s225  (
	.I0(\top/processor/sha_core/w[14] [12]),
	.I1(\top/processor/sha_core/w[15] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_139 )
);
defparam \top/processor/sha_core/n346_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s226  (
	.I0(\top/processor/sha_core/w[16] [12]),
	.I1(\top/processor/sha_core/w[17] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_140 )
);
defparam \top/processor/sha_core/n346_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s227  (
	.I0(\top/processor/sha_core/w[18] [12]),
	.I1(\top/processor/sha_core/w[19] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_141 )
);
defparam \top/processor/sha_core/n346_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s228  (
	.I0(\top/processor/sha_core/w[20] [12]),
	.I1(\top/processor/sha_core/w[21] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_142 )
);
defparam \top/processor/sha_core/n346_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s229  (
	.I0(\top/processor/sha_core/w[22] [12]),
	.I1(\top/processor/sha_core/w[23] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_143 )
);
defparam \top/processor/sha_core/n346_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s230  (
	.I0(\top/processor/sha_core/w[24] [12]),
	.I1(\top/processor/sha_core/w[25] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_144 )
);
defparam \top/processor/sha_core/n346_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s231  (
	.I0(\top/processor/sha_core/w[26] [12]),
	.I1(\top/processor/sha_core/w[27] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_145 )
);
defparam \top/processor/sha_core/n346_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s232  (
	.I0(\top/processor/sha_core/w[28] [12]),
	.I1(\top/processor/sha_core/w[29] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_146 )
);
defparam \top/processor/sha_core/n346_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s233  (
	.I0(\top/processor/sha_core/w[30] [12]),
	.I1(\top/processor/sha_core/w[31] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_147 )
);
defparam \top/processor/sha_core/n346_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s234  (
	.I0(\top/processor/sha_core/w[32] [12]),
	.I1(\top/processor/sha_core/w[33] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_148 )
);
defparam \top/processor/sha_core/n346_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s235  (
	.I0(\top/processor/sha_core/w[34] [12]),
	.I1(\top/processor/sha_core/w[35] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_149 )
);
defparam \top/processor/sha_core/n346_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s236  (
	.I0(\top/processor/sha_core/w[36] [12]),
	.I1(\top/processor/sha_core/w[37] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_150 )
);
defparam \top/processor/sha_core/n346_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s237  (
	.I0(\top/processor/sha_core/w[38] [12]),
	.I1(\top/processor/sha_core/w[39] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_151 )
);
defparam \top/processor/sha_core/n346_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s238  (
	.I0(\top/processor/sha_core/w[40] [12]),
	.I1(\top/processor/sha_core/w[41] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_152 )
);
defparam \top/processor/sha_core/n346_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s239  (
	.I0(\top/processor/sha_core/w[42] [12]),
	.I1(\top/processor/sha_core/w[43] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_153 )
);
defparam \top/processor/sha_core/n346_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s240  (
	.I0(\top/processor/sha_core/w[44] [12]),
	.I1(\top/processor/sha_core/w[45] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_154 )
);
defparam \top/processor/sha_core/n346_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s241  (
	.I0(\top/processor/sha_core/w[46] [12]),
	.I1(\top/processor/sha_core/w[47] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_155 )
);
defparam \top/processor/sha_core/n346_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s242  (
	.I0(\top/processor/sha_core/w[48] [12]),
	.I1(\top/processor/sha_core/w[49] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_156 )
);
defparam \top/processor/sha_core/n346_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s243  (
	.I0(\top/processor/sha_core/w[50] [12]),
	.I1(\top/processor/sha_core/w[51] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_157 )
);
defparam \top/processor/sha_core/n346_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s244  (
	.I0(\top/processor/sha_core/w[52] [12]),
	.I1(\top/processor/sha_core/w[53] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_158 )
);
defparam \top/processor/sha_core/n346_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s245  (
	.I0(\top/processor/sha_core/w[54] [12]),
	.I1(\top/processor/sha_core/w[55] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_159 )
);
defparam \top/processor/sha_core/n346_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s246  (
	.I0(\top/processor/sha_core/w[56] [12]),
	.I1(\top/processor/sha_core/w[57] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_160 )
);
defparam \top/processor/sha_core/n346_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s247  (
	.I0(\top/processor/sha_core/w[58] [12]),
	.I1(\top/processor/sha_core/w[59] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_161 )
);
defparam \top/processor/sha_core/n346_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s248  (
	.I0(\top/processor/sha_core/w[60] [12]),
	.I1(\top/processor/sha_core/w[61] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_162 )
);
defparam \top/processor/sha_core/n346_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s249  (
	.I0(\top/processor/sha_core/w[62] [12]),
	.I1(\top/processor/sha_core/w[63] [12]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n346_163 )
);
defparam \top/processor/sha_core/n346_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s218  (
	.I0(\top/processor/sha_core/w[0] [11]),
	.I1(\top/processor/sha_core/w[1] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_132 )
);
defparam \top/processor/sha_core/n347_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s219  (
	.I0(\top/processor/sha_core/w[2] [11]),
	.I1(\top/processor/sha_core/w[3] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_133 )
);
defparam \top/processor/sha_core/n347_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s220  (
	.I0(\top/processor/sha_core/w[4] [11]),
	.I1(\top/processor/sha_core/w[5] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_134 )
);
defparam \top/processor/sha_core/n347_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s221  (
	.I0(\top/processor/sha_core/w[6] [11]),
	.I1(\top/processor/sha_core/w[7] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_135 )
);
defparam \top/processor/sha_core/n347_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s222  (
	.I0(\top/processor/sha_core/w[8] [11]),
	.I1(\top/processor/sha_core/w[9] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_136 )
);
defparam \top/processor/sha_core/n347_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s223  (
	.I0(\top/processor/sha_core/w[10] [11]),
	.I1(\top/processor/sha_core/w[11] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_137 )
);
defparam \top/processor/sha_core/n347_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s224  (
	.I0(\top/processor/sha_core/w[12] [11]),
	.I1(\top/processor/sha_core/w[13] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_138 )
);
defparam \top/processor/sha_core/n347_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s225  (
	.I0(\top/processor/sha_core/w[14] [11]),
	.I1(\top/processor/sha_core/w[15] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_139 )
);
defparam \top/processor/sha_core/n347_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s226  (
	.I0(\top/processor/sha_core/w[16] [11]),
	.I1(\top/processor/sha_core/w[17] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_140 )
);
defparam \top/processor/sha_core/n347_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s227  (
	.I0(\top/processor/sha_core/w[18] [11]),
	.I1(\top/processor/sha_core/w[19] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_141 )
);
defparam \top/processor/sha_core/n347_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s228  (
	.I0(\top/processor/sha_core/w[20] [11]),
	.I1(\top/processor/sha_core/w[21] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_142 )
);
defparam \top/processor/sha_core/n347_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s229  (
	.I0(\top/processor/sha_core/w[22] [11]),
	.I1(\top/processor/sha_core/w[23] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_143 )
);
defparam \top/processor/sha_core/n347_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s230  (
	.I0(\top/processor/sha_core/w[24] [11]),
	.I1(\top/processor/sha_core/w[25] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_144 )
);
defparam \top/processor/sha_core/n347_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s231  (
	.I0(\top/processor/sha_core/w[26] [11]),
	.I1(\top/processor/sha_core/w[27] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_145 )
);
defparam \top/processor/sha_core/n347_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s232  (
	.I0(\top/processor/sha_core/w[28] [11]),
	.I1(\top/processor/sha_core/w[29] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_146 )
);
defparam \top/processor/sha_core/n347_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s233  (
	.I0(\top/processor/sha_core/w[30] [11]),
	.I1(\top/processor/sha_core/w[31] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_147 )
);
defparam \top/processor/sha_core/n347_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s234  (
	.I0(\top/processor/sha_core/w[32] [11]),
	.I1(\top/processor/sha_core/w[33] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_148 )
);
defparam \top/processor/sha_core/n347_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s235  (
	.I0(\top/processor/sha_core/w[34] [11]),
	.I1(\top/processor/sha_core/w[35] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_149 )
);
defparam \top/processor/sha_core/n347_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s236  (
	.I0(\top/processor/sha_core/w[36] [11]),
	.I1(\top/processor/sha_core/w[37] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_150 )
);
defparam \top/processor/sha_core/n347_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s237  (
	.I0(\top/processor/sha_core/w[38] [11]),
	.I1(\top/processor/sha_core/w[39] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_151 )
);
defparam \top/processor/sha_core/n347_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s238  (
	.I0(\top/processor/sha_core/w[40] [11]),
	.I1(\top/processor/sha_core/w[41] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_152 )
);
defparam \top/processor/sha_core/n347_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s239  (
	.I0(\top/processor/sha_core/w[42] [11]),
	.I1(\top/processor/sha_core/w[43] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_153 )
);
defparam \top/processor/sha_core/n347_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s240  (
	.I0(\top/processor/sha_core/w[44] [11]),
	.I1(\top/processor/sha_core/w[45] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_154 )
);
defparam \top/processor/sha_core/n347_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s241  (
	.I0(\top/processor/sha_core/w[46] [11]),
	.I1(\top/processor/sha_core/w[47] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_155 )
);
defparam \top/processor/sha_core/n347_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s242  (
	.I0(\top/processor/sha_core/w[48] [11]),
	.I1(\top/processor/sha_core/w[49] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_156 )
);
defparam \top/processor/sha_core/n347_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s243  (
	.I0(\top/processor/sha_core/w[50] [11]),
	.I1(\top/processor/sha_core/w[51] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_157 )
);
defparam \top/processor/sha_core/n347_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s244  (
	.I0(\top/processor/sha_core/w[52] [11]),
	.I1(\top/processor/sha_core/w[53] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_158 )
);
defparam \top/processor/sha_core/n347_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s245  (
	.I0(\top/processor/sha_core/w[54] [11]),
	.I1(\top/processor/sha_core/w[55] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_159 )
);
defparam \top/processor/sha_core/n347_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s246  (
	.I0(\top/processor/sha_core/w[56] [11]),
	.I1(\top/processor/sha_core/w[57] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_160 )
);
defparam \top/processor/sha_core/n347_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s247  (
	.I0(\top/processor/sha_core/w[58] [11]),
	.I1(\top/processor/sha_core/w[59] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_161 )
);
defparam \top/processor/sha_core/n347_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s248  (
	.I0(\top/processor/sha_core/w[60] [11]),
	.I1(\top/processor/sha_core/w[61] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_162 )
);
defparam \top/processor/sha_core/n347_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s249  (
	.I0(\top/processor/sha_core/w[62] [11]),
	.I1(\top/processor/sha_core/w[63] [11]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n347_163 )
);
defparam \top/processor/sha_core/n347_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s218  (
	.I0(\top/processor/sha_core/w[0] [10]),
	.I1(\top/processor/sha_core/w[1] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_132 )
);
defparam \top/processor/sha_core/n348_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s219  (
	.I0(\top/processor/sha_core/w[2] [10]),
	.I1(\top/processor/sha_core/w[3] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_133 )
);
defparam \top/processor/sha_core/n348_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s220  (
	.I0(\top/processor/sha_core/w[4] [10]),
	.I1(\top/processor/sha_core/w[5] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_134 )
);
defparam \top/processor/sha_core/n348_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s221  (
	.I0(\top/processor/sha_core/w[6] [10]),
	.I1(\top/processor/sha_core/w[7] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_135 )
);
defparam \top/processor/sha_core/n348_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s222  (
	.I0(\top/processor/sha_core/w[8] [10]),
	.I1(\top/processor/sha_core/w[9] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_136 )
);
defparam \top/processor/sha_core/n348_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s223  (
	.I0(\top/processor/sha_core/w[10] [10]),
	.I1(\top/processor/sha_core/w[11] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_137 )
);
defparam \top/processor/sha_core/n348_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s224  (
	.I0(\top/processor/sha_core/w[12] [10]),
	.I1(\top/processor/sha_core/w[13] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_138 )
);
defparam \top/processor/sha_core/n348_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s225  (
	.I0(\top/processor/sha_core/w[14] [10]),
	.I1(\top/processor/sha_core/w[15] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_139 )
);
defparam \top/processor/sha_core/n348_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s226  (
	.I0(\top/processor/sha_core/w[16] [10]),
	.I1(\top/processor/sha_core/w[17] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_140 )
);
defparam \top/processor/sha_core/n348_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s227  (
	.I0(\top/processor/sha_core/w[18] [10]),
	.I1(\top/processor/sha_core/w[19] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_141 )
);
defparam \top/processor/sha_core/n348_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s228  (
	.I0(\top/processor/sha_core/w[20] [10]),
	.I1(\top/processor/sha_core/w[21] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_142 )
);
defparam \top/processor/sha_core/n348_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s229  (
	.I0(\top/processor/sha_core/w[22] [10]),
	.I1(\top/processor/sha_core/w[23] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_143 )
);
defparam \top/processor/sha_core/n348_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s230  (
	.I0(\top/processor/sha_core/w[24] [10]),
	.I1(\top/processor/sha_core/w[25] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_144 )
);
defparam \top/processor/sha_core/n348_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s231  (
	.I0(\top/processor/sha_core/w[26] [10]),
	.I1(\top/processor/sha_core/w[27] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_145 )
);
defparam \top/processor/sha_core/n348_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s232  (
	.I0(\top/processor/sha_core/w[28] [10]),
	.I1(\top/processor/sha_core/w[29] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_146 )
);
defparam \top/processor/sha_core/n348_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s233  (
	.I0(\top/processor/sha_core/w[30] [10]),
	.I1(\top/processor/sha_core/w[31] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_147 )
);
defparam \top/processor/sha_core/n348_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s234  (
	.I0(\top/processor/sha_core/w[32] [10]),
	.I1(\top/processor/sha_core/w[33] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_148 )
);
defparam \top/processor/sha_core/n348_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s235  (
	.I0(\top/processor/sha_core/w[34] [10]),
	.I1(\top/processor/sha_core/w[35] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_149 )
);
defparam \top/processor/sha_core/n348_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s236  (
	.I0(\top/processor/sha_core/w[36] [10]),
	.I1(\top/processor/sha_core/w[37] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_150 )
);
defparam \top/processor/sha_core/n348_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s237  (
	.I0(\top/processor/sha_core/w[38] [10]),
	.I1(\top/processor/sha_core/w[39] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_151 )
);
defparam \top/processor/sha_core/n348_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s238  (
	.I0(\top/processor/sha_core/w[40] [10]),
	.I1(\top/processor/sha_core/w[41] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_152 )
);
defparam \top/processor/sha_core/n348_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s239  (
	.I0(\top/processor/sha_core/w[42] [10]),
	.I1(\top/processor/sha_core/w[43] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_153 )
);
defparam \top/processor/sha_core/n348_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s240  (
	.I0(\top/processor/sha_core/w[44] [10]),
	.I1(\top/processor/sha_core/w[45] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_154 )
);
defparam \top/processor/sha_core/n348_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s241  (
	.I0(\top/processor/sha_core/w[46] [10]),
	.I1(\top/processor/sha_core/w[47] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_155 )
);
defparam \top/processor/sha_core/n348_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s242  (
	.I0(\top/processor/sha_core/w[48] [10]),
	.I1(\top/processor/sha_core/w[49] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_156 )
);
defparam \top/processor/sha_core/n348_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s243  (
	.I0(\top/processor/sha_core/w[50] [10]),
	.I1(\top/processor/sha_core/w[51] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_157 )
);
defparam \top/processor/sha_core/n348_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s244  (
	.I0(\top/processor/sha_core/w[52] [10]),
	.I1(\top/processor/sha_core/w[53] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_158 )
);
defparam \top/processor/sha_core/n348_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s245  (
	.I0(\top/processor/sha_core/w[54] [10]),
	.I1(\top/processor/sha_core/w[55] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_159 )
);
defparam \top/processor/sha_core/n348_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s246  (
	.I0(\top/processor/sha_core/w[56] [10]),
	.I1(\top/processor/sha_core/w[57] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_160 )
);
defparam \top/processor/sha_core/n348_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s247  (
	.I0(\top/processor/sha_core/w[58] [10]),
	.I1(\top/processor/sha_core/w[59] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_161 )
);
defparam \top/processor/sha_core/n348_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s248  (
	.I0(\top/processor/sha_core/w[60] [10]),
	.I1(\top/processor/sha_core/w[61] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_162 )
);
defparam \top/processor/sha_core/n348_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s249  (
	.I0(\top/processor/sha_core/w[62] [10]),
	.I1(\top/processor/sha_core/w[63] [10]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n348_163 )
);
defparam \top/processor/sha_core/n348_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s218  (
	.I0(\top/processor/sha_core/w[0] [9]),
	.I1(\top/processor/sha_core/w[1] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_132 )
);
defparam \top/processor/sha_core/n349_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s219  (
	.I0(\top/processor/sha_core/w[2] [9]),
	.I1(\top/processor/sha_core/w[3] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_133 )
);
defparam \top/processor/sha_core/n349_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s220  (
	.I0(\top/processor/sha_core/w[4] [9]),
	.I1(\top/processor/sha_core/w[5] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_134 )
);
defparam \top/processor/sha_core/n349_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s221  (
	.I0(\top/processor/sha_core/w[6] [9]),
	.I1(\top/processor/sha_core/w[7] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_135 )
);
defparam \top/processor/sha_core/n349_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s222  (
	.I0(\top/processor/sha_core/w[8] [9]),
	.I1(\top/processor/sha_core/w[9] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_136 )
);
defparam \top/processor/sha_core/n349_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s223  (
	.I0(\top/processor/sha_core/w[10] [9]),
	.I1(\top/processor/sha_core/w[11] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_137 )
);
defparam \top/processor/sha_core/n349_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s224  (
	.I0(\top/processor/sha_core/w[12] [9]),
	.I1(\top/processor/sha_core/w[13] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_138 )
);
defparam \top/processor/sha_core/n349_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s225  (
	.I0(\top/processor/sha_core/w[14] [9]),
	.I1(\top/processor/sha_core/w[15] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_139 )
);
defparam \top/processor/sha_core/n349_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s226  (
	.I0(\top/processor/sha_core/w[16] [9]),
	.I1(\top/processor/sha_core/w[17] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_140 )
);
defparam \top/processor/sha_core/n349_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s227  (
	.I0(\top/processor/sha_core/w[18] [9]),
	.I1(\top/processor/sha_core/w[19] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_141 )
);
defparam \top/processor/sha_core/n349_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s228  (
	.I0(\top/processor/sha_core/w[20] [9]),
	.I1(\top/processor/sha_core/w[21] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_142 )
);
defparam \top/processor/sha_core/n349_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s229  (
	.I0(\top/processor/sha_core/w[22] [9]),
	.I1(\top/processor/sha_core/w[23] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_143 )
);
defparam \top/processor/sha_core/n349_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s230  (
	.I0(\top/processor/sha_core/w[24] [9]),
	.I1(\top/processor/sha_core/w[25] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_144 )
);
defparam \top/processor/sha_core/n349_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s231  (
	.I0(\top/processor/sha_core/w[26] [9]),
	.I1(\top/processor/sha_core/w[27] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_145 )
);
defparam \top/processor/sha_core/n349_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s232  (
	.I0(\top/processor/sha_core/w[28] [9]),
	.I1(\top/processor/sha_core/w[29] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_146 )
);
defparam \top/processor/sha_core/n349_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s233  (
	.I0(\top/processor/sha_core/w[30] [9]),
	.I1(\top/processor/sha_core/w[31] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_147 )
);
defparam \top/processor/sha_core/n349_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s234  (
	.I0(\top/processor/sha_core/w[32] [9]),
	.I1(\top/processor/sha_core/w[33] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_148 )
);
defparam \top/processor/sha_core/n349_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s235  (
	.I0(\top/processor/sha_core/w[34] [9]),
	.I1(\top/processor/sha_core/w[35] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_149 )
);
defparam \top/processor/sha_core/n349_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s236  (
	.I0(\top/processor/sha_core/w[36] [9]),
	.I1(\top/processor/sha_core/w[37] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_150 )
);
defparam \top/processor/sha_core/n349_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s237  (
	.I0(\top/processor/sha_core/w[38] [9]),
	.I1(\top/processor/sha_core/w[39] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_151 )
);
defparam \top/processor/sha_core/n349_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s238  (
	.I0(\top/processor/sha_core/w[40] [9]),
	.I1(\top/processor/sha_core/w[41] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_152 )
);
defparam \top/processor/sha_core/n349_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s239  (
	.I0(\top/processor/sha_core/w[42] [9]),
	.I1(\top/processor/sha_core/w[43] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_153 )
);
defparam \top/processor/sha_core/n349_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s240  (
	.I0(\top/processor/sha_core/w[44] [9]),
	.I1(\top/processor/sha_core/w[45] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_154 )
);
defparam \top/processor/sha_core/n349_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s241  (
	.I0(\top/processor/sha_core/w[46] [9]),
	.I1(\top/processor/sha_core/w[47] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_155 )
);
defparam \top/processor/sha_core/n349_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s242  (
	.I0(\top/processor/sha_core/w[48] [9]),
	.I1(\top/processor/sha_core/w[49] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_156 )
);
defparam \top/processor/sha_core/n349_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s243  (
	.I0(\top/processor/sha_core/w[50] [9]),
	.I1(\top/processor/sha_core/w[51] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_157 )
);
defparam \top/processor/sha_core/n349_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s244  (
	.I0(\top/processor/sha_core/w[52] [9]),
	.I1(\top/processor/sha_core/w[53] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_158 )
);
defparam \top/processor/sha_core/n349_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s245  (
	.I0(\top/processor/sha_core/w[54] [9]),
	.I1(\top/processor/sha_core/w[55] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_159 )
);
defparam \top/processor/sha_core/n349_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s246  (
	.I0(\top/processor/sha_core/w[56] [9]),
	.I1(\top/processor/sha_core/w[57] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_160 )
);
defparam \top/processor/sha_core/n349_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s247  (
	.I0(\top/processor/sha_core/w[58] [9]),
	.I1(\top/processor/sha_core/w[59] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_161 )
);
defparam \top/processor/sha_core/n349_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s248  (
	.I0(\top/processor/sha_core/w[60] [9]),
	.I1(\top/processor/sha_core/w[61] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_162 )
);
defparam \top/processor/sha_core/n349_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s249  (
	.I0(\top/processor/sha_core/w[62] [9]),
	.I1(\top/processor/sha_core/w[63] [9]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n349_163 )
);
defparam \top/processor/sha_core/n349_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s218  (
	.I0(\top/processor/sha_core/w[0] [8]),
	.I1(\top/processor/sha_core/w[1] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_132 )
);
defparam \top/processor/sha_core/n350_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s219  (
	.I0(\top/processor/sha_core/w[2] [8]),
	.I1(\top/processor/sha_core/w[3] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_133 )
);
defparam \top/processor/sha_core/n350_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s220  (
	.I0(\top/processor/sha_core/w[4] [8]),
	.I1(\top/processor/sha_core/w[5] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_134 )
);
defparam \top/processor/sha_core/n350_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s221  (
	.I0(\top/processor/sha_core/w[6] [8]),
	.I1(\top/processor/sha_core/w[7] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_135 )
);
defparam \top/processor/sha_core/n350_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s222  (
	.I0(\top/processor/sha_core/w[8] [8]),
	.I1(\top/processor/sha_core/w[9] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_136 )
);
defparam \top/processor/sha_core/n350_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s223  (
	.I0(\top/processor/sha_core/w[10] [8]),
	.I1(\top/processor/sha_core/w[11] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_137 )
);
defparam \top/processor/sha_core/n350_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s224  (
	.I0(\top/processor/sha_core/w[12] [8]),
	.I1(\top/processor/sha_core/w[13] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_138 )
);
defparam \top/processor/sha_core/n350_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s225  (
	.I0(\top/processor/sha_core/w[14] [8]),
	.I1(\top/processor/sha_core/w[15] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_139 )
);
defparam \top/processor/sha_core/n350_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s226  (
	.I0(\top/processor/sha_core/w[16] [8]),
	.I1(\top/processor/sha_core/w[17] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_140 )
);
defparam \top/processor/sha_core/n350_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s227  (
	.I0(\top/processor/sha_core/w[18] [8]),
	.I1(\top/processor/sha_core/w[19] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_141 )
);
defparam \top/processor/sha_core/n350_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s228  (
	.I0(\top/processor/sha_core/w[20] [8]),
	.I1(\top/processor/sha_core/w[21] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_142 )
);
defparam \top/processor/sha_core/n350_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s229  (
	.I0(\top/processor/sha_core/w[22] [8]),
	.I1(\top/processor/sha_core/w[23] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_143 )
);
defparam \top/processor/sha_core/n350_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s230  (
	.I0(\top/processor/sha_core/w[24] [8]),
	.I1(\top/processor/sha_core/w[25] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_144 )
);
defparam \top/processor/sha_core/n350_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s231  (
	.I0(\top/processor/sha_core/w[26] [8]),
	.I1(\top/processor/sha_core/w[27] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_145 )
);
defparam \top/processor/sha_core/n350_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s232  (
	.I0(\top/processor/sha_core/w[28] [8]),
	.I1(\top/processor/sha_core/w[29] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_146 )
);
defparam \top/processor/sha_core/n350_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s233  (
	.I0(\top/processor/sha_core/w[30] [8]),
	.I1(\top/processor/sha_core/w[31] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_147 )
);
defparam \top/processor/sha_core/n350_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s234  (
	.I0(\top/processor/sha_core/w[32] [8]),
	.I1(\top/processor/sha_core/w[33] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_148 )
);
defparam \top/processor/sha_core/n350_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s235  (
	.I0(\top/processor/sha_core/w[34] [8]),
	.I1(\top/processor/sha_core/w[35] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_149 )
);
defparam \top/processor/sha_core/n350_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s236  (
	.I0(\top/processor/sha_core/w[36] [8]),
	.I1(\top/processor/sha_core/w[37] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_150 )
);
defparam \top/processor/sha_core/n350_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s237  (
	.I0(\top/processor/sha_core/w[38] [8]),
	.I1(\top/processor/sha_core/w[39] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_151 )
);
defparam \top/processor/sha_core/n350_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s238  (
	.I0(\top/processor/sha_core/w[40] [8]),
	.I1(\top/processor/sha_core/w[41] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_152 )
);
defparam \top/processor/sha_core/n350_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s239  (
	.I0(\top/processor/sha_core/w[42] [8]),
	.I1(\top/processor/sha_core/w[43] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_153 )
);
defparam \top/processor/sha_core/n350_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s240  (
	.I0(\top/processor/sha_core/w[44] [8]),
	.I1(\top/processor/sha_core/w[45] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_154 )
);
defparam \top/processor/sha_core/n350_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s241  (
	.I0(\top/processor/sha_core/w[46] [8]),
	.I1(\top/processor/sha_core/w[47] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_155 )
);
defparam \top/processor/sha_core/n350_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s242  (
	.I0(\top/processor/sha_core/w[48] [8]),
	.I1(\top/processor/sha_core/w[49] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_156 )
);
defparam \top/processor/sha_core/n350_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s243  (
	.I0(\top/processor/sha_core/w[50] [8]),
	.I1(\top/processor/sha_core/w[51] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_157 )
);
defparam \top/processor/sha_core/n350_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s244  (
	.I0(\top/processor/sha_core/w[52] [8]),
	.I1(\top/processor/sha_core/w[53] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_158 )
);
defparam \top/processor/sha_core/n350_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s245  (
	.I0(\top/processor/sha_core/w[54] [8]),
	.I1(\top/processor/sha_core/w[55] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_159 )
);
defparam \top/processor/sha_core/n350_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s246  (
	.I0(\top/processor/sha_core/w[56] [8]),
	.I1(\top/processor/sha_core/w[57] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_160 )
);
defparam \top/processor/sha_core/n350_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s247  (
	.I0(\top/processor/sha_core/w[58] [8]),
	.I1(\top/processor/sha_core/w[59] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_161 )
);
defparam \top/processor/sha_core/n350_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s248  (
	.I0(\top/processor/sha_core/w[60] [8]),
	.I1(\top/processor/sha_core/w[61] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_162 )
);
defparam \top/processor/sha_core/n350_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s249  (
	.I0(\top/processor/sha_core/w[62] [8]),
	.I1(\top/processor/sha_core/w[63] [8]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n350_163 )
);
defparam \top/processor/sha_core/n350_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s218  (
	.I0(\top/processor/sha_core/w[0] [7]),
	.I1(\top/processor/sha_core/w[1] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_132 )
);
defparam \top/processor/sha_core/n351_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s219  (
	.I0(\top/processor/sha_core/w[2] [7]),
	.I1(\top/processor/sha_core/w[3] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_133 )
);
defparam \top/processor/sha_core/n351_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s220  (
	.I0(\top/processor/sha_core/w[4] [7]),
	.I1(\top/processor/sha_core/w[5] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_134 )
);
defparam \top/processor/sha_core/n351_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s221  (
	.I0(\top/processor/sha_core/w[6] [7]),
	.I1(\top/processor/sha_core/w[7] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_135 )
);
defparam \top/processor/sha_core/n351_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s222  (
	.I0(\top/processor/sha_core/w[8] [7]),
	.I1(\top/processor/sha_core/w[9] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_136 )
);
defparam \top/processor/sha_core/n351_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s223  (
	.I0(\top/processor/sha_core/w[10] [7]),
	.I1(\top/processor/sha_core/w[11] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_137 )
);
defparam \top/processor/sha_core/n351_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s224  (
	.I0(\top/processor/sha_core/w[12] [7]),
	.I1(\top/processor/sha_core/w[13] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_138 )
);
defparam \top/processor/sha_core/n351_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s225  (
	.I0(\top/processor/sha_core/w[14] [7]),
	.I1(\top/processor/sha_core/w[15] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_139 )
);
defparam \top/processor/sha_core/n351_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s226  (
	.I0(\top/processor/sha_core/w[16] [7]),
	.I1(\top/processor/sha_core/w[17] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_140 )
);
defparam \top/processor/sha_core/n351_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s227  (
	.I0(\top/processor/sha_core/w[18] [7]),
	.I1(\top/processor/sha_core/w[19] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_141 )
);
defparam \top/processor/sha_core/n351_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s228  (
	.I0(\top/processor/sha_core/w[20] [7]),
	.I1(\top/processor/sha_core/w[21] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_142 )
);
defparam \top/processor/sha_core/n351_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s229  (
	.I0(\top/processor/sha_core/w[22] [7]),
	.I1(\top/processor/sha_core/w[23] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_143 )
);
defparam \top/processor/sha_core/n351_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s230  (
	.I0(\top/processor/sha_core/w[24] [7]),
	.I1(\top/processor/sha_core/w[25] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_144 )
);
defparam \top/processor/sha_core/n351_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s231  (
	.I0(\top/processor/sha_core/w[26] [7]),
	.I1(\top/processor/sha_core/w[27] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_145 )
);
defparam \top/processor/sha_core/n351_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s232  (
	.I0(\top/processor/sha_core/w[28] [7]),
	.I1(\top/processor/sha_core/w[29] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_146 )
);
defparam \top/processor/sha_core/n351_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s233  (
	.I0(\top/processor/sha_core/w[30] [7]),
	.I1(\top/processor/sha_core/w[31] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_147 )
);
defparam \top/processor/sha_core/n351_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s234  (
	.I0(\top/processor/sha_core/w[32] [7]),
	.I1(\top/processor/sha_core/w[33] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_148 )
);
defparam \top/processor/sha_core/n351_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s235  (
	.I0(\top/processor/sha_core/w[34] [7]),
	.I1(\top/processor/sha_core/w[35] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_149 )
);
defparam \top/processor/sha_core/n351_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s236  (
	.I0(\top/processor/sha_core/w[36] [7]),
	.I1(\top/processor/sha_core/w[37] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_150 )
);
defparam \top/processor/sha_core/n351_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s237  (
	.I0(\top/processor/sha_core/w[38] [7]),
	.I1(\top/processor/sha_core/w[39] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_151 )
);
defparam \top/processor/sha_core/n351_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s238  (
	.I0(\top/processor/sha_core/w[40] [7]),
	.I1(\top/processor/sha_core/w[41] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_152 )
);
defparam \top/processor/sha_core/n351_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s239  (
	.I0(\top/processor/sha_core/w[42] [7]),
	.I1(\top/processor/sha_core/w[43] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_153 )
);
defparam \top/processor/sha_core/n351_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s240  (
	.I0(\top/processor/sha_core/w[44] [7]),
	.I1(\top/processor/sha_core/w[45] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_154 )
);
defparam \top/processor/sha_core/n351_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s241  (
	.I0(\top/processor/sha_core/w[46] [7]),
	.I1(\top/processor/sha_core/w[47] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_155 )
);
defparam \top/processor/sha_core/n351_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s242  (
	.I0(\top/processor/sha_core/w[48] [7]),
	.I1(\top/processor/sha_core/w[49] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_156 )
);
defparam \top/processor/sha_core/n351_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s243  (
	.I0(\top/processor/sha_core/w[50] [7]),
	.I1(\top/processor/sha_core/w[51] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_157 )
);
defparam \top/processor/sha_core/n351_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s244  (
	.I0(\top/processor/sha_core/w[52] [7]),
	.I1(\top/processor/sha_core/w[53] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_158 )
);
defparam \top/processor/sha_core/n351_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s245  (
	.I0(\top/processor/sha_core/w[54] [7]),
	.I1(\top/processor/sha_core/w[55] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_159 )
);
defparam \top/processor/sha_core/n351_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s246  (
	.I0(\top/processor/sha_core/w[56] [7]),
	.I1(\top/processor/sha_core/w[57] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_160 )
);
defparam \top/processor/sha_core/n351_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s247  (
	.I0(\top/processor/sha_core/w[58] [7]),
	.I1(\top/processor/sha_core/w[59] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_161 )
);
defparam \top/processor/sha_core/n351_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s248  (
	.I0(\top/processor/sha_core/w[60] [7]),
	.I1(\top/processor/sha_core/w[61] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_162 )
);
defparam \top/processor/sha_core/n351_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s249  (
	.I0(\top/processor/sha_core/w[62] [7]),
	.I1(\top/processor/sha_core/w[63] [7]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n351_163 )
);
defparam \top/processor/sha_core/n351_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s218  (
	.I0(\top/processor/sha_core/w[0] [6]),
	.I1(\top/processor/sha_core/w[1] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_132 )
);
defparam \top/processor/sha_core/n352_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s219  (
	.I0(\top/processor/sha_core/w[2] [6]),
	.I1(\top/processor/sha_core/w[3] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_133 )
);
defparam \top/processor/sha_core/n352_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s220  (
	.I0(\top/processor/sha_core/w[4] [6]),
	.I1(\top/processor/sha_core/w[5] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_134 )
);
defparam \top/processor/sha_core/n352_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s221  (
	.I0(\top/processor/sha_core/w[6] [6]),
	.I1(\top/processor/sha_core/w[7] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_135 )
);
defparam \top/processor/sha_core/n352_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s222  (
	.I0(\top/processor/sha_core/w[8] [6]),
	.I1(\top/processor/sha_core/w[9] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_136 )
);
defparam \top/processor/sha_core/n352_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s223  (
	.I0(\top/processor/sha_core/w[10] [6]),
	.I1(\top/processor/sha_core/w[11] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_137 )
);
defparam \top/processor/sha_core/n352_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s224  (
	.I0(\top/processor/sha_core/w[12] [6]),
	.I1(\top/processor/sha_core/w[13] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_138 )
);
defparam \top/processor/sha_core/n352_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s225  (
	.I0(\top/processor/sha_core/w[14] [6]),
	.I1(\top/processor/sha_core/w[15] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_139 )
);
defparam \top/processor/sha_core/n352_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s226  (
	.I0(\top/processor/sha_core/w[16] [6]),
	.I1(\top/processor/sha_core/w[17] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_140 )
);
defparam \top/processor/sha_core/n352_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s227  (
	.I0(\top/processor/sha_core/w[18] [6]),
	.I1(\top/processor/sha_core/w[19] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_141 )
);
defparam \top/processor/sha_core/n352_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s228  (
	.I0(\top/processor/sha_core/w[20] [6]),
	.I1(\top/processor/sha_core/w[21] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_142 )
);
defparam \top/processor/sha_core/n352_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s229  (
	.I0(\top/processor/sha_core/w[22] [6]),
	.I1(\top/processor/sha_core/w[23] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_143 )
);
defparam \top/processor/sha_core/n352_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s230  (
	.I0(\top/processor/sha_core/w[24] [6]),
	.I1(\top/processor/sha_core/w[25] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_144 )
);
defparam \top/processor/sha_core/n352_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s231  (
	.I0(\top/processor/sha_core/w[26] [6]),
	.I1(\top/processor/sha_core/w[27] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_145 )
);
defparam \top/processor/sha_core/n352_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s232  (
	.I0(\top/processor/sha_core/w[28] [6]),
	.I1(\top/processor/sha_core/w[29] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_146 )
);
defparam \top/processor/sha_core/n352_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s233  (
	.I0(\top/processor/sha_core/w[30] [6]),
	.I1(\top/processor/sha_core/w[31] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_147 )
);
defparam \top/processor/sha_core/n352_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s234  (
	.I0(\top/processor/sha_core/w[32] [6]),
	.I1(\top/processor/sha_core/w[33] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_148 )
);
defparam \top/processor/sha_core/n352_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s235  (
	.I0(\top/processor/sha_core/w[34] [6]),
	.I1(\top/processor/sha_core/w[35] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_149 )
);
defparam \top/processor/sha_core/n352_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s236  (
	.I0(\top/processor/sha_core/w[36] [6]),
	.I1(\top/processor/sha_core/w[37] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_150 )
);
defparam \top/processor/sha_core/n352_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s237  (
	.I0(\top/processor/sha_core/w[38] [6]),
	.I1(\top/processor/sha_core/w[39] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_151 )
);
defparam \top/processor/sha_core/n352_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s238  (
	.I0(\top/processor/sha_core/w[40] [6]),
	.I1(\top/processor/sha_core/w[41] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_152 )
);
defparam \top/processor/sha_core/n352_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s239  (
	.I0(\top/processor/sha_core/w[42] [6]),
	.I1(\top/processor/sha_core/w[43] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_153 )
);
defparam \top/processor/sha_core/n352_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s240  (
	.I0(\top/processor/sha_core/w[44] [6]),
	.I1(\top/processor/sha_core/w[45] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_154 )
);
defparam \top/processor/sha_core/n352_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s241  (
	.I0(\top/processor/sha_core/w[46] [6]),
	.I1(\top/processor/sha_core/w[47] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_155 )
);
defparam \top/processor/sha_core/n352_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s242  (
	.I0(\top/processor/sha_core/w[48] [6]),
	.I1(\top/processor/sha_core/w[49] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_156 )
);
defparam \top/processor/sha_core/n352_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s243  (
	.I0(\top/processor/sha_core/w[50] [6]),
	.I1(\top/processor/sha_core/w[51] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_157 )
);
defparam \top/processor/sha_core/n352_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s244  (
	.I0(\top/processor/sha_core/w[52] [6]),
	.I1(\top/processor/sha_core/w[53] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_158 )
);
defparam \top/processor/sha_core/n352_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s245  (
	.I0(\top/processor/sha_core/w[54] [6]),
	.I1(\top/processor/sha_core/w[55] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_159 )
);
defparam \top/processor/sha_core/n352_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s246  (
	.I0(\top/processor/sha_core/w[56] [6]),
	.I1(\top/processor/sha_core/w[57] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_160 )
);
defparam \top/processor/sha_core/n352_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s247  (
	.I0(\top/processor/sha_core/w[58] [6]),
	.I1(\top/processor/sha_core/w[59] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_161 )
);
defparam \top/processor/sha_core/n352_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s248  (
	.I0(\top/processor/sha_core/w[60] [6]),
	.I1(\top/processor/sha_core/w[61] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_162 )
);
defparam \top/processor/sha_core/n352_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s249  (
	.I0(\top/processor/sha_core/w[62] [6]),
	.I1(\top/processor/sha_core/w[63] [6]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n352_163 )
);
defparam \top/processor/sha_core/n352_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s218  (
	.I0(\top/processor/sha_core/w[0] [5]),
	.I1(\top/processor/sha_core/w[1] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_132 )
);
defparam \top/processor/sha_core/n353_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s219  (
	.I0(\top/processor/sha_core/w[2] [5]),
	.I1(\top/processor/sha_core/w[3] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_133 )
);
defparam \top/processor/sha_core/n353_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s220  (
	.I0(\top/processor/sha_core/w[4] [5]),
	.I1(\top/processor/sha_core/w[5] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_134 )
);
defparam \top/processor/sha_core/n353_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s221  (
	.I0(\top/processor/sha_core/w[6] [5]),
	.I1(\top/processor/sha_core/w[7] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_135 )
);
defparam \top/processor/sha_core/n353_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s222  (
	.I0(\top/processor/sha_core/w[8] [5]),
	.I1(\top/processor/sha_core/w[9] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_136 )
);
defparam \top/processor/sha_core/n353_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s223  (
	.I0(\top/processor/sha_core/w[10] [5]),
	.I1(\top/processor/sha_core/w[11] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_137 )
);
defparam \top/processor/sha_core/n353_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s224  (
	.I0(\top/processor/sha_core/w[12] [5]),
	.I1(\top/processor/sha_core/w[13] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_138 )
);
defparam \top/processor/sha_core/n353_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s225  (
	.I0(\top/processor/sha_core/w[14] [5]),
	.I1(\top/processor/sha_core/w[15] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_139 )
);
defparam \top/processor/sha_core/n353_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s226  (
	.I0(\top/processor/sha_core/w[16] [5]),
	.I1(\top/processor/sha_core/w[17] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_140 )
);
defparam \top/processor/sha_core/n353_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s227  (
	.I0(\top/processor/sha_core/w[18] [5]),
	.I1(\top/processor/sha_core/w[19] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_141 )
);
defparam \top/processor/sha_core/n353_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s228  (
	.I0(\top/processor/sha_core/w[20] [5]),
	.I1(\top/processor/sha_core/w[21] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_142 )
);
defparam \top/processor/sha_core/n353_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s229  (
	.I0(\top/processor/sha_core/w[22] [5]),
	.I1(\top/processor/sha_core/w[23] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_143 )
);
defparam \top/processor/sha_core/n353_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s230  (
	.I0(\top/processor/sha_core/w[24] [5]),
	.I1(\top/processor/sha_core/w[25] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_144 )
);
defparam \top/processor/sha_core/n353_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s231  (
	.I0(\top/processor/sha_core/w[26] [5]),
	.I1(\top/processor/sha_core/w[27] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_145 )
);
defparam \top/processor/sha_core/n353_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s232  (
	.I0(\top/processor/sha_core/w[28] [5]),
	.I1(\top/processor/sha_core/w[29] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_146 )
);
defparam \top/processor/sha_core/n353_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s233  (
	.I0(\top/processor/sha_core/w[30] [5]),
	.I1(\top/processor/sha_core/w[31] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_147 )
);
defparam \top/processor/sha_core/n353_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s234  (
	.I0(\top/processor/sha_core/w[32] [5]),
	.I1(\top/processor/sha_core/w[33] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_148 )
);
defparam \top/processor/sha_core/n353_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s235  (
	.I0(\top/processor/sha_core/w[34] [5]),
	.I1(\top/processor/sha_core/w[35] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_149 )
);
defparam \top/processor/sha_core/n353_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s236  (
	.I0(\top/processor/sha_core/w[36] [5]),
	.I1(\top/processor/sha_core/w[37] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_150 )
);
defparam \top/processor/sha_core/n353_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s237  (
	.I0(\top/processor/sha_core/w[38] [5]),
	.I1(\top/processor/sha_core/w[39] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_151 )
);
defparam \top/processor/sha_core/n353_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s238  (
	.I0(\top/processor/sha_core/w[40] [5]),
	.I1(\top/processor/sha_core/w[41] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_152 )
);
defparam \top/processor/sha_core/n353_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s239  (
	.I0(\top/processor/sha_core/w[42] [5]),
	.I1(\top/processor/sha_core/w[43] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_153 )
);
defparam \top/processor/sha_core/n353_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s240  (
	.I0(\top/processor/sha_core/w[44] [5]),
	.I1(\top/processor/sha_core/w[45] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_154 )
);
defparam \top/processor/sha_core/n353_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s241  (
	.I0(\top/processor/sha_core/w[46] [5]),
	.I1(\top/processor/sha_core/w[47] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_155 )
);
defparam \top/processor/sha_core/n353_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s242  (
	.I0(\top/processor/sha_core/w[48] [5]),
	.I1(\top/processor/sha_core/w[49] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_156 )
);
defparam \top/processor/sha_core/n353_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s243  (
	.I0(\top/processor/sha_core/w[50] [5]),
	.I1(\top/processor/sha_core/w[51] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_157 )
);
defparam \top/processor/sha_core/n353_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s244  (
	.I0(\top/processor/sha_core/w[52] [5]),
	.I1(\top/processor/sha_core/w[53] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_158 )
);
defparam \top/processor/sha_core/n353_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s245  (
	.I0(\top/processor/sha_core/w[54] [5]),
	.I1(\top/processor/sha_core/w[55] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_159 )
);
defparam \top/processor/sha_core/n353_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s246  (
	.I0(\top/processor/sha_core/w[56] [5]),
	.I1(\top/processor/sha_core/w[57] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_160 )
);
defparam \top/processor/sha_core/n353_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s247  (
	.I0(\top/processor/sha_core/w[58] [5]),
	.I1(\top/processor/sha_core/w[59] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_161 )
);
defparam \top/processor/sha_core/n353_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s248  (
	.I0(\top/processor/sha_core/w[60] [5]),
	.I1(\top/processor/sha_core/w[61] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_162 )
);
defparam \top/processor/sha_core/n353_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s249  (
	.I0(\top/processor/sha_core/w[62] [5]),
	.I1(\top/processor/sha_core/w[63] [5]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n353_163 )
);
defparam \top/processor/sha_core/n353_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s218  (
	.I0(\top/processor/sha_core/w[0] [4]),
	.I1(\top/processor/sha_core/w[1] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_132 )
);
defparam \top/processor/sha_core/n354_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s219  (
	.I0(\top/processor/sha_core/w[2] [4]),
	.I1(\top/processor/sha_core/w[3] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_133 )
);
defparam \top/processor/sha_core/n354_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s220  (
	.I0(\top/processor/sha_core/w[4] [4]),
	.I1(\top/processor/sha_core/w[5] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_134 )
);
defparam \top/processor/sha_core/n354_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s221  (
	.I0(\top/processor/sha_core/w[6] [4]),
	.I1(\top/processor/sha_core/w[7] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_135 )
);
defparam \top/processor/sha_core/n354_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s222  (
	.I0(\top/processor/sha_core/w[8] [4]),
	.I1(\top/processor/sha_core/w[9] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_136 )
);
defparam \top/processor/sha_core/n354_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s223  (
	.I0(\top/processor/sha_core/w[10] [4]),
	.I1(\top/processor/sha_core/w[11] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_137 )
);
defparam \top/processor/sha_core/n354_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s224  (
	.I0(\top/processor/sha_core/w[12] [4]),
	.I1(\top/processor/sha_core/w[13] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_138 )
);
defparam \top/processor/sha_core/n354_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s225  (
	.I0(\top/processor/sha_core/w[14] [4]),
	.I1(\top/processor/sha_core/w[15] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_139 )
);
defparam \top/processor/sha_core/n354_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s226  (
	.I0(\top/processor/sha_core/w[16] [4]),
	.I1(\top/processor/sha_core/w[17] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_140 )
);
defparam \top/processor/sha_core/n354_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s227  (
	.I0(\top/processor/sha_core/w[18] [4]),
	.I1(\top/processor/sha_core/w[19] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_141 )
);
defparam \top/processor/sha_core/n354_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s228  (
	.I0(\top/processor/sha_core/w[20] [4]),
	.I1(\top/processor/sha_core/w[21] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_142 )
);
defparam \top/processor/sha_core/n354_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s229  (
	.I0(\top/processor/sha_core/w[22] [4]),
	.I1(\top/processor/sha_core/w[23] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_143 )
);
defparam \top/processor/sha_core/n354_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s230  (
	.I0(\top/processor/sha_core/w[24] [4]),
	.I1(\top/processor/sha_core/w[25] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_144 )
);
defparam \top/processor/sha_core/n354_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s231  (
	.I0(\top/processor/sha_core/w[26] [4]),
	.I1(\top/processor/sha_core/w[27] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_145 )
);
defparam \top/processor/sha_core/n354_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s232  (
	.I0(\top/processor/sha_core/w[28] [4]),
	.I1(\top/processor/sha_core/w[29] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_146 )
);
defparam \top/processor/sha_core/n354_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s233  (
	.I0(\top/processor/sha_core/w[30] [4]),
	.I1(\top/processor/sha_core/w[31] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_147 )
);
defparam \top/processor/sha_core/n354_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s234  (
	.I0(\top/processor/sha_core/w[32] [4]),
	.I1(\top/processor/sha_core/w[33] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_148 )
);
defparam \top/processor/sha_core/n354_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s235  (
	.I0(\top/processor/sha_core/w[34] [4]),
	.I1(\top/processor/sha_core/w[35] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_149 )
);
defparam \top/processor/sha_core/n354_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s236  (
	.I0(\top/processor/sha_core/w[36] [4]),
	.I1(\top/processor/sha_core/w[37] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_150 )
);
defparam \top/processor/sha_core/n354_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s237  (
	.I0(\top/processor/sha_core/w[38] [4]),
	.I1(\top/processor/sha_core/w[39] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_151 )
);
defparam \top/processor/sha_core/n354_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s238  (
	.I0(\top/processor/sha_core/w[40] [4]),
	.I1(\top/processor/sha_core/w[41] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_152 )
);
defparam \top/processor/sha_core/n354_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s239  (
	.I0(\top/processor/sha_core/w[42] [4]),
	.I1(\top/processor/sha_core/w[43] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_153 )
);
defparam \top/processor/sha_core/n354_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s240  (
	.I0(\top/processor/sha_core/w[44] [4]),
	.I1(\top/processor/sha_core/w[45] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_154 )
);
defparam \top/processor/sha_core/n354_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s241  (
	.I0(\top/processor/sha_core/w[46] [4]),
	.I1(\top/processor/sha_core/w[47] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_155 )
);
defparam \top/processor/sha_core/n354_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s242  (
	.I0(\top/processor/sha_core/w[48] [4]),
	.I1(\top/processor/sha_core/w[49] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_156 )
);
defparam \top/processor/sha_core/n354_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s243  (
	.I0(\top/processor/sha_core/w[50] [4]),
	.I1(\top/processor/sha_core/w[51] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_157 )
);
defparam \top/processor/sha_core/n354_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s244  (
	.I0(\top/processor/sha_core/w[52] [4]),
	.I1(\top/processor/sha_core/w[53] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_158 )
);
defparam \top/processor/sha_core/n354_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s245  (
	.I0(\top/processor/sha_core/w[54] [4]),
	.I1(\top/processor/sha_core/w[55] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_159 )
);
defparam \top/processor/sha_core/n354_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s246  (
	.I0(\top/processor/sha_core/w[56] [4]),
	.I1(\top/processor/sha_core/w[57] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_160 )
);
defparam \top/processor/sha_core/n354_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s247  (
	.I0(\top/processor/sha_core/w[58] [4]),
	.I1(\top/processor/sha_core/w[59] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_161 )
);
defparam \top/processor/sha_core/n354_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s248  (
	.I0(\top/processor/sha_core/w[60] [4]),
	.I1(\top/processor/sha_core/w[61] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_162 )
);
defparam \top/processor/sha_core/n354_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s249  (
	.I0(\top/processor/sha_core/w[62] [4]),
	.I1(\top/processor/sha_core/w[63] [4]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n354_163 )
);
defparam \top/processor/sha_core/n354_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s218  (
	.I0(\top/processor/sha_core/w[0] [3]),
	.I1(\top/processor/sha_core/w[1] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_132 )
);
defparam \top/processor/sha_core/n355_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s219  (
	.I0(\top/processor/sha_core/w[2] [3]),
	.I1(\top/processor/sha_core/w[3] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_133 )
);
defparam \top/processor/sha_core/n355_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s220  (
	.I0(\top/processor/sha_core/w[4] [3]),
	.I1(\top/processor/sha_core/w[5] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_134 )
);
defparam \top/processor/sha_core/n355_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s221  (
	.I0(\top/processor/sha_core/w[6] [3]),
	.I1(\top/processor/sha_core/w[7] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_135 )
);
defparam \top/processor/sha_core/n355_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s222  (
	.I0(\top/processor/sha_core/w[8] [3]),
	.I1(\top/processor/sha_core/w[9] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_136 )
);
defparam \top/processor/sha_core/n355_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s223  (
	.I0(\top/processor/sha_core/w[10] [3]),
	.I1(\top/processor/sha_core/w[11] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_137 )
);
defparam \top/processor/sha_core/n355_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s224  (
	.I0(\top/processor/sha_core/w[12] [3]),
	.I1(\top/processor/sha_core/w[13] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_138 )
);
defparam \top/processor/sha_core/n355_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s225  (
	.I0(\top/processor/sha_core/w[14] [3]),
	.I1(\top/processor/sha_core/w[15] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_139 )
);
defparam \top/processor/sha_core/n355_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s226  (
	.I0(\top/processor/sha_core/w[16] [3]),
	.I1(\top/processor/sha_core/w[17] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_140 )
);
defparam \top/processor/sha_core/n355_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s227  (
	.I0(\top/processor/sha_core/w[18] [3]),
	.I1(\top/processor/sha_core/w[19] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_141 )
);
defparam \top/processor/sha_core/n355_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s228  (
	.I0(\top/processor/sha_core/w[20] [3]),
	.I1(\top/processor/sha_core/w[21] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_142 )
);
defparam \top/processor/sha_core/n355_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s229  (
	.I0(\top/processor/sha_core/w[22] [3]),
	.I1(\top/processor/sha_core/w[23] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_143 )
);
defparam \top/processor/sha_core/n355_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s230  (
	.I0(\top/processor/sha_core/w[24] [3]),
	.I1(\top/processor/sha_core/w[25] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_144 )
);
defparam \top/processor/sha_core/n355_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s231  (
	.I0(\top/processor/sha_core/w[26] [3]),
	.I1(\top/processor/sha_core/w[27] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_145 )
);
defparam \top/processor/sha_core/n355_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s232  (
	.I0(\top/processor/sha_core/w[28] [3]),
	.I1(\top/processor/sha_core/w[29] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_146 )
);
defparam \top/processor/sha_core/n355_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s233  (
	.I0(\top/processor/sha_core/w[30] [3]),
	.I1(\top/processor/sha_core/w[31] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_147 )
);
defparam \top/processor/sha_core/n355_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s234  (
	.I0(\top/processor/sha_core/w[32] [3]),
	.I1(\top/processor/sha_core/w[33] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_148 )
);
defparam \top/processor/sha_core/n355_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s235  (
	.I0(\top/processor/sha_core/w[34] [3]),
	.I1(\top/processor/sha_core/w[35] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_149 )
);
defparam \top/processor/sha_core/n355_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s236  (
	.I0(\top/processor/sha_core/w[36] [3]),
	.I1(\top/processor/sha_core/w[37] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_150 )
);
defparam \top/processor/sha_core/n355_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s237  (
	.I0(\top/processor/sha_core/w[38] [3]),
	.I1(\top/processor/sha_core/w[39] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_151 )
);
defparam \top/processor/sha_core/n355_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s238  (
	.I0(\top/processor/sha_core/w[40] [3]),
	.I1(\top/processor/sha_core/w[41] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_152 )
);
defparam \top/processor/sha_core/n355_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s239  (
	.I0(\top/processor/sha_core/w[42] [3]),
	.I1(\top/processor/sha_core/w[43] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_153 )
);
defparam \top/processor/sha_core/n355_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s240  (
	.I0(\top/processor/sha_core/w[44] [3]),
	.I1(\top/processor/sha_core/w[45] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_154 )
);
defparam \top/processor/sha_core/n355_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s241  (
	.I0(\top/processor/sha_core/w[46] [3]),
	.I1(\top/processor/sha_core/w[47] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_155 )
);
defparam \top/processor/sha_core/n355_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s242  (
	.I0(\top/processor/sha_core/w[48] [3]),
	.I1(\top/processor/sha_core/w[49] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_156 )
);
defparam \top/processor/sha_core/n355_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s243  (
	.I0(\top/processor/sha_core/w[50] [3]),
	.I1(\top/processor/sha_core/w[51] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_157 )
);
defparam \top/processor/sha_core/n355_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s244  (
	.I0(\top/processor/sha_core/w[52] [3]),
	.I1(\top/processor/sha_core/w[53] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_158 )
);
defparam \top/processor/sha_core/n355_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s245  (
	.I0(\top/processor/sha_core/w[54] [3]),
	.I1(\top/processor/sha_core/w[55] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_159 )
);
defparam \top/processor/sha_core/n355_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s246  (
	.I0(\top/processor/sha_core/w[56] [3]),
	.I1(\top/processor/sha_core/w[57] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_160 )
);
defparam \top/processor/sha_core/n355_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s247  (
	.I0(\top/processor/sha_core/w[58] [3]),
	.I1(\top/processor/sha_core/w[59] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_161 )
);
defparam \top/processor/sha_core/n355_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s248  (
	.I0(\top/processor/sha_core/w[60] [3]),
	.I1(\top/processor/sha_core/w[61] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_162 )
);
defparam \top/processor/sha_core/n355_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s249  (
	.I0(\top/processor/sha_core/w[62] [3]),
	.I1(\top/processor/sha_core/w[63] [3]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n355_163 )
);
defparam \top/processor/sha_core/n355_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s218  (
	.I0(\top/processor/sha_core/w[0] [2]),
	.I1(\top/processor/sha_core/w[1] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_132 )
);
defparam \top/processor/sha_core/n356_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s219  (
	.I0(\top/processor/sha_core/w[2] [2]),
	.I1(\top/processor/sha_core/w[3] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_133 )
);
defparam \top/processor/sha_core/n356_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s220  (
	.I0(\top/processor/sha_core/w[4] [2]),
	.I1(\top/processor/sha_core/w[5] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_134 )
);
defparam \top/processor/sha_core/n356_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s221  (
	.I0(\top/processor/sha_core/w[6] [2]),
	.I1(\top/processor/sha_core/w[7] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_135 )
);
defparam \top/processor/sha_core/n356_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s222  (
	.I0(\top/processor/sha_core/w[8] [2]),
	.I1(\top/processor/sha_core/w[9] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_136 )
);
defparam \top/processor/sha_core/n356_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s223  (
	.I0(\top/processor/sha_core/w[10] [2]),
	.I1(\top/processor/sha_core/w[11] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_137 )
);
defparam \top/processor/sha_core/n356_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s224  (
	.I0(\top/processor/sha_core/w[12] [2]),
	.I1(\top/processor/sha_core/w[13] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_138 )
);
defparam \top/processor/sha_core/n356_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s225  (
	.I0(\top/processor/sha_core/w[14] [2]),
	.I1(\top/processor/sha_core/w[15] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_139 )
);
defparam \top/processor/sha_core/n356_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s226  (
	.I0(\top/processor/sha_core/w[16] [2]),
	.I1(\top/processor/sha_core/w[17] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_140 )
);
defparam \top/processor/sha_core/n356_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s227  (
	.I0(\top/processor/sha_core/w[18] [2]),
	.I1(\top/processor/sha_core/w[19] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_141 )
);
defparam \top/processor/sha_core/n356_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s228  (
	.I0(\top/processor/sha_core/w[20] [2]),
	.I1(\top/processor/sha_core/w[21] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_142 )
);
defparam \top/processor/sha_core/n356_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s229  (
	.I0(\top/processor/sha_core/w[22] [2]),
	.I1(\top/processor/sha_core/w[23] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_143 )
);
defparam \top/processor/sha_core/n356_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s230  (
	.I0(\top/processor/sha_core/w[24] [2]),
	.I1(\top/processor/sha_core/w[25] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_144 )
);
defparam \top/processor/sha_core/n356_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s231  (
	.I0(\top/processor/sha_core/w[26] [2]),
	.I1(\top/processor/sha_core/w[27] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_145 )
);
defparam \top/processor/sha_core/n356_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s232  (
	.I0(\top/processor/sha_core/w[28] [2]),
	.I1(\top/processor/sha_core/w[29] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_146 )
);
defparam \top/processor/sha_core/n356_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s233  (
	.I0(\top/processor/sha_core/w[30] [2]),
	.I1(\top/processor/sha_core/w[31] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_147 )
);
defparam \top/processor/sha_core/n356_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s234  (
	.I0(\top/processor/sha_core/w[32] [2]),
	.I1(\top/processor/sha_core/w[33] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_148 )
);
defparam \top/processor/sha_core/n356_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s235  (
	.I0(\top/processor/sha_core/w[34] [2]),
	.I1(\top/processor/sha_core/w[35] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_149 )
);
defparam \top/processor/sha_core/n356_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s236  (
	.I0(\top/processor/sha_core/w[36] [2]),
	.I1(\top/processor/sha_core/w[37] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_150 )
);
defparam \top/processor/sha_core/n356_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s237  (
	.I0(\top/processor/sha_core/w[38] [2]),
	.I1(\top/processor/sha_core/w[39] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_151 )
);
defparam \top/processor/sha_core/n356_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s238  (
	.I0(\top/processor/sha_core/w[40] [2]),
	.I1(\top/processor/sha_core/w[41] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_152 )
);
defparam \top/processor/sha_core/n356_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s239  (
	.I0(\top/processor/sha_core/w[42] [2]),
	.I1(\top/processor/sha_core/w[43] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_153 )
);
defparam \top/processor/sha_core/n356_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s240  (
	.I0(\top/processor/sha_core/w[44] [2]),
	.I1(\top/processor/sha_core/w[45] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_154 )
);
defparam \top/processor/sha_core/n356_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s241  (
	.I0(\top/processor/sha_core/w[46] [2]),
	.I1(\top/processor/sha_core/w[47] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_155 )
);
defparam \top/processor/sha_core/n356_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s242  (
	.I0(\top/processor/sha_core/w[48] [2]),
	.I1(\top/processor/sha_core/w[49] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_156 )
);
defparam \top/processor/sha_core/n356_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s243  (
	.I0(\top/processor/sha_core/w[50] [2]),
	.I1(\top/processor/sha_core/w[51] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_157 )
);
defparam \top/processor/sha_core/n356_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s244  (
	.I0(\top/processor/sha_core/w[52] [2]),
	.I1(\top/processor/sha_core/w[53] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_158 )
);
defparam \top/processor/sha_core/n356_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s245  (
	.I0(\top/processor/sha_core/w[54] [2]),
	.I1(\top/processor/sha_core/w[55] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_159 )
);
defparam \top/processor/sha_core/n356_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s246  (
	.I0(\top/processor/sha_core/w[56] [2]),
	.I1(\top/processor/sha_core/w[57] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_160 )
);
defparam \top/processor/sha_core/n356_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s247  (
	.I0(\top/processor/sha_core/w[58] [2]),
	.I1(\top/processor/sha_core/w[59] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_161 )
);
defparam \top/processor/sha_core/n356_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s248  (
	.I0(\top/processor/sha_core/w[60] [2]),
	.I1(\top/processor/sha_core/w[61] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_162 )
);
defparam \top/processor/sha_core/n356_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s249  (
	.I0(\top/processor/sha_core/w[62] [2]),
	.I1(\top/processor/sha_core/w[63] [2]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n356_163 )
);
defparam \top/processor/sha_core/n356_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s218  (
	.I0(\top/processor/sha_core/w[0] [1]),
	.I1(\top/processor/sha_core/w[1] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_132 )
);
defparam \top/processor/sha_core/n357_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s219  (
	.I0(\top/processor/sha_core/w[2] [1]),
	.I1(\top/processor/sha_core/w[3] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_133 )
);
defparam \top/processor/sha_core/n357_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s220  (
	.I0(\top/processor/sha_core/w[4] [1]),
	.I1(\top/processor/sha_core/w[5] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_134 )
);
defparam \top/processor/sha_core/n357_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s221  (
	.I0(\top/processor/sha_core/w[6] [1]),
	.I1(\top/processor/sha_core/w[7] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_135 )
);
defparam \top/processor/sha_core/n357_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s222  (
	.I0(\top/processor/sha_core/w[8] [1]),
	.I1(\top/processor/sha_core/w[9] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_136 )
);
defparam \top/processor/sha_core/n357_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s223  (
	.I0(\top/processor/sha_core/w[10] [1]),
	.I1(\top/processor/sha_core/w[11] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_137 )
);
defparam \top/processor/sha_core/n357_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s224  (
	.I0(\top/processor/sha_core/w[12] [1]),
	.I1(\top/processor/sha_core/w[13] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_138 )
);
defparam \top/processor/sha_core/n357_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s225  (
	.I0(\top/processor/sha_core/w[14] [1]),
	.I1(\top/processor/sha_core/w[15] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_139 )
);
defparam \top/processor/sha_core/n357_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s226  (
	.I0(\top/processor/sha_core/w[16] [1]),
	.I1(\top/processor/sha_core/w[17] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_140 )
);
defparam \top/processor/sha_core/n357_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s227  (
	.I0(\top/processor/sha_core/w[18] [1]),
	.I1(\top/processor/sha_core/w[19] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_141 )
);
defparam \top/processor/sha_core/n357_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s228  (
	.I0(\top/processor/sha_core/w[20] [1]),
	.I1(\top/processor/sha_core/w[21] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_142 )
);
defparam \top/processor/sha_core/n357_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s229  (
	.I0(\top/processor/sha_core/w[22] [1]),
	.I1(\top/processor/sha_core/w[23] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_143 )
);
defparam \top/processor/sha_core/n357_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s230  (
	.I0(\top/processor/sha_core/w[24] [1]),
	.I1(\top/processor/sha_core/w[25] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_144 )
);
defparam \top/processor/sha_core/n357_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s231  (
	.I0(\top/processor/sha_core/w[26] [1]),
	.I1(\top/processor/sha_core/w[27] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_145 )
);
defparam \top/processor/sha_core/n357_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s232  (
	.I0(\top/processor/sha_core/w[28] [1]),
	.I1(\top/processor/sha_core/w[29] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_146 )
);
defparam \top/processor/sha_core/n357_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s233  (
	.I0(\top/processor/sha_core/w[30] [1]),
	.I1(\top/processor/sha_core/w[31] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_147 )
);
defparam \top/processor/sha_core/n357_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s234  (
	.I0(\top/processor/sha_core/w[32] [1]),
	.I1(\top/processor/sha_core/w[33] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_148 )
);
defparam \top/processor/sha_core/n357_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s235  (
	.I0(\top/processor/sha_core/w[34] [1]),
	.I1(\top/processor/sha_core/w[35] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_149 )
);
defparam \top/processor/sha_core/n357_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s236  (
	.I0(\top/processor/sha_core/w[36] [1]),
	.I1(\top/processor/sha_core/w[37] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_150 )
);
defparam \top/processor/sha_core/n357_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s237  (
	.I0(\top/processor/sha_core/w[38] [1]),
	.I1(\top/processor/sha_core/w[39] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_151 )
);
defparam \top/processor/sha_core/n357_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s238  (
	.I0(\top/processor/sha_core/w[40] [1]),
	.I1(\top/processor/sha_core/w[41] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_152 )
);
defparam \top/processor/sha_core/n357_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s239  (
	.I0(\top/processor/sha_core/w[42] [1]),
	.I1(\top/processor/sha_core/w[43] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_153 )
);
defparam \top/processor/sha_core/n357_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s240  (
	.I0(\top/processor/sha_core/w[44] [1]),
	.I1(\top/processor/sha_core/w[45] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_154 )
);
defparam \top/processor/sha_core/n357_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s241  (
	.I0(\top/processor/sha_core/w[46] [1]),
	.I1(\top/processor/sha_core/w[47] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_155 )
);
defparam \top/processor/sha_core/n357_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s242  (
	.I0(\top/processor/sha_core/w[48] [1]),
	.I1(\top/processor/sha_core/w[49] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_156 )
);
defparam \top/processor/sha_core/n357_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s243  (
	.I0(\top/processor/sha_core/w[50] [1]),
	.I1(\top/processor/sha_core/w[51] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_157 )
);
defparam \top/processor/sha_core/n357_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s244  (
	.I0(\top/processor/sha_core/w[52] [1]),
	.I1(\top/processor/sha_core/w[53] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_158 )
);
defparam \top/processor/sha_core/n357_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s245  (
	.I0(\top/processor/sha_core/w[54] [1]),
	.I1(\top/processor/sha_core/w[55] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_159 )
);
defparam \top/processor/sha_core/n357_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s246  (
	.I0(\top/processor/sha_core/w[56] [1]),
	.I1(\top/processor/sha_core/w[57] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_160 )
);
defparam \top/processor/sha_core/n357_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s247  (
	.I0(\top/processor/sha_core/w[58] [1]),
	.I1(\top/processor/sha_core/w[59] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_161 )
);
defparam \top/processor/sha_core/n357_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s248  (
	.I0(\top/processor/sha_core/w[60] [1]),
	.I1(\top/processor/sha_core/w[61] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_162 )
);
defparam \top/processor/sha_core/n357_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s249  (
	.I0(\top/processor/sha_core/w[62] [1]),
	.I1(\top/processor/sha_core/w[63] [1]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n357_163 )
);
defparam \top/processor/sha_core/n357_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s218  (
	.I0(\top/processor/sha_core/w[0] [0]),
	.I1(\top/processor/sha_core/w[1] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_132 )
);
defparam \top/processor/sha_core/n358_s218 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s219  (
	.I0(\top/processor/sha_core/w[2] [0]),
	.I1(\top/processor/sha_core/w[3] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_133 )
);
defparam \top/processor/sha_core/n358_s219 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s220  (
	.I0(\top/processor/sha_core/w[4] [0]),
	.I1(\top/processor/sha_core/w[5] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_134 )
);
defparam \top/processor/sha_core/n358_s220 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s221  (
	.I0(\top/processor/sha_core/w[6] [0]),
	.I1(\top/processor/sha_core/w[7] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_135 )
);
defparam \top/processor/sha_core/n358_s221 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s222  (
	.I0(\top/processor/sha_core/w[8] [0]),
	.I1(\top/processor/sha_core/w[9] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_136 )
);
defparam \top/processor/sha_core/n358_s222 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s223  (
	.I0(\top/processor/sha_core/w[10] [0]),
	.I1(\top/processor/sha_core/w[11] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_137 )
);
defparam \top/processor/sha_core/n358_s223 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s224  (
	.I0(\top/processor/sha_core/w[12] [0]),
	.I1(\top/processor/sha_core/w[13] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_138 )
);
defparam \top/processor/sha_core/n358_s224 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s225  (
	.I0(\top/processor/sha_core/w[14] [0]),
	.I1(\top/processor/sha_core/w[15] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_139 )
);
defparam \top/processor/sha_core/n358_s225 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s226  (
	.I0(\top/processor/sha_core/w[16] [0]),
	.I1(\top/processor/sha_core/w[17] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_140 )
);
defparam \top/processor/sha_core/n358_s226 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s227  (
	.I0(\top/processor/sha_core/w[18] [0]),
	.I1(\top/processor/sha_core/w[19] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_141 )
);
defparam \top/processor/sha_core/n358_s227 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s228  (
	.I0(\top/processor/sha_core/w[20] [0]),
	.I1(\top/processor/sha_core/w[21] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_142 )
);
defparam \top/processor/sha_core/n358_s228 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s229  (
	.I0(\top/processor/sha_core/w[22] [0]),
	.I1(\top/processor/sha_core/w[23] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_143 )
);
defparam \top/processor/sha_core/n358_s229 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s230  (
	.I0(\top/processor/sha_core/w[24] [0]),
	.I1(\top/processor/sha_core/w[25] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_144 )
);
defparam \top/processor/sha_core/n358_s230 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s231  (
	.I0(\top/processor/sha_core/w[26] [0]),
	.I1(\top/processor/sha_core/w[27] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_145 )
);
defparam \top/processor/sha_core/n358_s231 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s232  (
	.I0(\top/processor/sha_core/w[28] [0]),
	.I1(\top/processor/sha_core/w[29] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_146 )
);
defparam \top/processor/sha_core/n358_s232 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s233  (
	.I0(\top/processor/sha_core/w[30] [0]),
	.I1(\top/processor/sha_core/w[31] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_147 )
);
defparam \top/processor/sha_core/n358_s233 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s234  (
	.I0(\top/processor/sha_core/w[32] [0]),
	.I1(\top/processor/sha_core/w[33] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_148 )
);
defparam \top/processor/sha_core/n358_s234 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s235  (
	.I0(\top/processor/sha_core/w[34] [0]),
	.I1(\top/processor/sha_core/w[35] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_149 )
);
defparam \top/processor/sha_core/n358_s235 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s236  (
	.I0(\top/processor/sha_core/w[36] [0]),
	.I1(\top/processor/sha_core/w[37] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_150 )
);
defparam \top/processor/sha_core/n358_s236 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s237  (
	.I0(\top/processor/sha_core/w[38] [0]),
	.I1(\top/processor/sha_core/w[39] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_151 )
);
defparam \top/processor/sha_core/n358_s237 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s238  (
	.I0(\top/processor/sha_core/w[40] [0]),
	.I1(\top/processor/sha_core/w[41] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_152 )
);
defparam \top/processor/sha_core/n358_s238 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s239  (
	.I0(\top/processor/sha_core/w[42] [0]),
	.I1(\top/processor/sha_core/w[43] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_153 )
);
defparam \top/processor/sha_core/n358_s239 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s240  (
	.I0(\top/processor/sha_core/w[44] [0]),
	.I1(\top/processor/sha_core/w[45] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_154 )
);
defparam \top/processor/sha_core/n358_s240 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s241  (
	.I0(\top/processor/sha_core/w[46] [0]),
	.I1(\top/processor/sha_core/w[47] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_155 )
);
defparam \top/processor/sha_core/n358_s241 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s242  (
	.I0(\top/processor/sha_core/w[48] [0]),
	.I1(\top/processor/sha_core/w[49] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_156 )
);
defparam \top/processor/sha_core/n358_s242 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s243  (
	.I0(\top/processor/sha_core/w[50] [0]),
	.I1(\top/processor/sha_core/w[51] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_157 )
);
defparam \top/processor/sha_core/n358_s243 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s244  (
	.I0(\top/processor/sha_core/w[52] [0]),
	.I1(\top/processor/sha_core/w[53] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_158 )
);
defparam \top/processor/sha_core/n358_s244 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s245  (
	.I0(\top/processor/sha_core/w[54] [0]),
	.I1(\top/processor/sha_core/w[55] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_159 )
);
defparam \top/processor/sha_core/n358_s245 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s246  (
	.I0(\top/processor/sha_core/w[56] [0]),
	.I1(\top/processor/sha_core/w[57] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_160 )
);
defparam \top/processor/sha_core/n358_s246 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s247  (
	.I0(\top/processor/sha_core/w[58] [0]),
	.I1(\top/processor/sha_core/w[59] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_161 )
);
defparam \top/processor/sha_core/n358_s247 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s248  (
	.I0(\top/processor/sha_core/w[60] [0]),
	.I1(\top/processor/sha_core/w[61] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_162 )
);
defparam \top/processor/sha_core/n358_s248 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s249  (
	.I0(\top/processor/sha_core/w[62] [0]),
	.I1(\top/processor/sha_core/w[63] [0]),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n358_163 )
);
defparam \top/processor/sha_core/n358_s249 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n36_s0  (
	.I0(\top/processor/sha_core/e [6]),
	.I1(\top/processor/sha_core/e [11]),
	.I2(\top/processor/sha_core/e [25]),
	.F(\top/processor/sha_core/n36_3 )
);
defparam \top/processor/sha_core/n36_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n37_s0  (
	.I0(\top/processor/sha_core/e [7]),
	.I1(\top/processor/sha_core/e [12]),
	.I2(\top/processor/sha_core/e [26]),
	.F(\top/processor/sha_core/n37_3 )
);
defparam \top/processor/sha_core/n37_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n38_s0  (
	.I0(\top/processor/sha_core/e [8]),
	.I1(\top/processor/sha_core/e [13]),
	.I2(\top/processor/sha_core/e [27]),
	.F(\top/processor/sha_core/n38_3 )
);
defparam \top/processor/sha_core/n38_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n39_s0  (
	.I0(\top/processor/sha_core/e [9]),
	.I1(\top/processor/sha_core/e [14]),
	.I2(\top/processor/sha_core/e [28]),
	.F(\top/processor/sha_core/n39_3 )
);
defparam \top/processor/sha_core/n39_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n40_s0  (
	.I0(\top/processor/sha_core/e [10]),
	.I1(\top/processor/sha_core/e [15]),
	.I2(\top/processor/sha_core/e [29]),
	.F(\top/processor/sha_core/n40_3 )
);
defparam \top/processor/sha_core/n40_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n41_s0  (
	.I0(\top/processor/sha_core/e [11]),
	.I1(\top/processor/sha_core/e [16]),
	.I2(\top/processor/sha_core/e [30]),
	.F(\top/processor/sha_core/n41_3 )
);
defparam \top/processor/sha_core/n41_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n42_s0  (
	.I0(\top/processor/sha_core/e [12]),
	.I1(\top/processor/sha_core/e [17]),
	.I2(\top/processor/sha_core/e [31]),
	.F(\top/processor/sha_core/n42_3 )
);
defparam \top/processor/sha_core/n42_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n43_s0  (
	.I0(\top/processor/sha_core/e [13]),
	.I1(\top/processor/sha_core/e [18]),
	.I2(\top/processor/sha_core/e [0]),
	.F(\top/processor/sha_core/n43_3 )
);
defparam \top/processor/sha_core/n43_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n44_s0  (
	.I0(\top/processor/sha_core/e [14]),
	.I1(\top/processor/sha_core/e [19]),
	.I2(\top/processor/sha_core/e [1]),
	.F(\top/processor/sha_core/n44_3 )
);
defparam \top/processor/sha_core/n44_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n45_s0  (
	.I0(\top/processor/sha_core/e [15]),
	.I1(\top/processor/sha_core/e [20]),
	.I2(\top/processor/sha_core/e [2]),
	.F(\top/processor/sha_core/n45_3 )
);
defparam \top/processor/sha_core/n45_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n46_s0  (
	.I0(\top/processor/sha_core/e [16]),
	.I1(\top/processor/sha_core/e [21]),
	.I2(\top/processor/sha_core/e [3]),
	.F(\top/processor/sha_core/n46_3 )
);
defparam \top/processor/sha_core/n46_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n47_s0  (
	.I0(\top/processor/sha_core/e [17]),
	.I1(\top/processor/sha_core/e [22]),
	.I2(\top/processor/sha_core/e [4]),
	.F(\top/processor/sha_core/n47_3 )
);
defparam \top/processor/sha_core/n47_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n48_s0  (
	.I0(\top/processor/sha_core/e [18]),
	.I1(\top/processor/sha_core/e [23]),
	.I2(\top/processor/sha_core/e [5]),
	.F(\top/processor/sha_core/n48_3 )
);
defparam \top/processor/sha_core/n48_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n49_s0  (
	.I0(\top/processor/sha_core/e [6]),
	.I1(\top/processor/sha_core/e [19]),
	.I2(\top/processor/sha_core/e [24]),
	.F(\top/processor/sha_core/n49_3 )
);
defparam \top/processor/sha_core/n49_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n50_s0  (
	.I0(\top/processor/sha_core/e [7]),
	.I1(\top/processor/sha_core/e [20]),
	.I2(\top/processor/sha_core/e [25]),
	.F(\top/processor/sha_core/n50_3 )
);
defparam \top/processor/sha_core/n50_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n51_s0  (
	.I0(\top/processor/sha_core/e [8]),
	.I1(\top/processor/sha_core/e [21]),
	.I2(\top/processor/sha_core/e [26]),
	.F(\top/processor/sha_core/n51_3 )
);
defparam \top/processor/sha_core/n51_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n52_s0  (
	.I0(\top/processor/sha_core/e [9]),
	.I1(\top/processor/sha_core/e [22]),
	.I2(\top/processor/sha_core/e [27]),
	.F(\top/processor/sha_core/n52_3 )
);
defparam \top/processor/sha_core/n52_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n53_s0  (
	.I0(\top/processor/sha_core/e [10]),
	.I1(\top/processor/sha_core/e [23]),
	.I2(\top/processor/sha_core/e [28]),
	.F(\top/processor/sha_core/n53_3 )
);
defparam \top/processor/sha_core/n53_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n54_s0  (
	.I0(\top/processor/sha_core/e [11]),
	.I1(\top/processor/sha_core/e [24]),
	.I2(\top/processor/sha_core/e [29]),
	.F(\top/processor/sha_core/n54_3 )
);
defparam \top/processor/sha_core/n54_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n55_s0  (
	.I0(\top/processor/sha_core/e [12]),
	.I1(\top/processor/sha_core/e [25]),
	.I2(\top/processor/sha_core/e [30]),
	.F(\top/processor/sha_core/n55_3 )
);
defparam \top/processor/sha_core/n55_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n56_s0  (
	.I0(\top/processor/sha_core/e [13]),
	.I1(\top/processor/sha_core/e [26]),
	.I2(\top/processor/sha_core/e [31]),
	.F(\top/processor/sha_core/n56_3 )
);
defparam \top/processor/sha_core/n56_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n57_s0  (
	.I0(\top/processor/sha_core/e [14]),
	.I1(\top/processor/sha_core/e [27]),
	.I2(\top/processor/sha_core/e [0]),
	.F(\top/processor/sha_core/n57_3 )
);
defparam \top/processor/sha_core/n57_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n58_s0  (
	.I0(\top/processor/sha_core/e [15]),
	.I1(\top/processor/sha_core/e [28]),
	.I2(\top/processor/sha_core/e [1]),
	.F(\top/processor/sha_core/n58_3 )
);
defparam \top/processor/sha_core/n58_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n59_s0  (
	.I0(\top/processor/sha_core/e [16]),
	.I1(\top/processor/sha_core/e [29]),
	.I2(\top/processor/sha_core/e [2]),
	.F(\top/processor/sha_core/n59_3 )
);
defparam \top/processor/sha_core/n59_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n60_s0  (
	.I0(\top/processor/sha_core/e [17]),
	.I1(\top/processor/sha_core/e [30]),
	.I2(\top/processor/sha_core/e [3]),
	.F(\top/processor/sha_core/n60_3 )
);
defparam \top/processor/sha_core/n60_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n61_s0  (
	.I0(\top/processor/sha_core/e [18]),
	.I1(\top/processor/sha_core/e [31]),
	.I2(\top/processor/sha_core/e [4]),
	.F(\top/processor/sha_core/n61_3 )
);
defparam \top/processor/sha_core/n61_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n62_s0  (
	.I0(\top/processor/sha_core/e [19]),
	.I1(\top/processor/sha_core/e [0]),
	.I2(\top/processor/sha_core/e [5]),
	.F(\top/processor/sha_core/n62_3 )
);
defparam \top/processor/sha_core/n62_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n63_s0  (
	.I0(\top/processor/sha_core/e [6]),
	.I1(\top/processor/sha_core/e [20]),
	.I2(\top/processor/sha_core/e [1]),
	.F(\top/processor/sha_core/n63_3 )
);
defparam \top/processor/sha_core/n63_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n64_s0  (
	.I0(\top/processor/sha_core/e [7]),
	.I1(\top/processor/sha_core/e [21]),
	.I2(\top/processor/sha_core/e [2]),
	.F(\top/processor/sha_core/n64_3 )
);
defparam \top/processor/sha_core/n64_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n65_s0  (
	.I0(\top/processor/sha_core/e [8]),
	.I1(\top/processor/sha_core/e [22]),
	.I2(\top/processor/sha_core/e [3]),
	.F(\top/processor/sha_core/n65_3 )
);
defparam \top/processor/sha_core/n65_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n66_s0  (
	.I0(\top/processor/sha_core/e [9]),
	.I1(\top/processor/sha_core/e [23]),
	.I2(\top/processor/sha_core/e [4]),
	.F(\top/processor/sha_core/n66_3 )
);
defparam \top/processor/sha_core/n66_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n67_s0  (
	.I0(\top/processor/sha_core/e [10]),
	.I1(\top/processor/sha_core/e [24]),
	.I2(\top/processor/sha_core/e [5]),
	.F(\top/processor/sha_core/n67_3 )
);
defparam \top/processor/sha_core/n67_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n197_s0  (
	.I0(\top/processor/sha_core/g [0]),
	.I1(\top/processor/sha_core/f [0]),
	.I2(\top/processor/sha_core/e [0]),
	.F(\top/processor/sha_core/n197_3 )
);
defparam \top/processor/sha_core/n197_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n198_s0  (
	.I0(\top/processor/sha_core/g [1]),
	.I1(\top/processor/sha_core/f [1]),
	.I2(\top/processor/sha_core/e [1]),
	.F(\top/processor/sha_core/n198_3 )
);
defparam \top/processor/sha_core/n198_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n199_s0  (
	.I0(\top/processor/sha_core/g [2]),
	.I1(\top/processor/sha_core/f [2]),
	.I2(\top/processor/sha_core/e [2]),
	.F(\top/processor/sha_core/n199_3 )
);
defparam \top/processor/sha_core/n199_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n200_s0  (
	.I0(\top/processor/sha_core/g [3]),
	.I1(\top/processor/sha_core/f [3]),
	.I2(\top/processor/sha_core/e [3]),
	.F(\top/processor/sha_core/n200_3 )
);
defparam \top/processor/sha_core/n200_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n201_s0  (
	.I0(\top/processor/sha_core/g [4]),
	.I1(\top/processor/sha_core/f [4]),
	.I2(\top/processor/sha_core/e [4]),
	.F(\top/processor/sha_core/n201_3 )
);
defparam \top/processor/sha_core/n201_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n202_s0  (
	.I0(\top/processor/sha_core/g [5]),
	.I1(\top/processor/sha_core/f [5]),
	.I2(\top/processor/sha_core/e [5]),
	.F(\top/processor/sha_core/n202_3 )
);
defparam \top/processor/sha_core/n202_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n203_s0  (
	.I0(\top/processor/sha_core/g [6]),
	.I1(\top/processor/sha_core/f [6]),
	.I2(\top/processor/sha_core/e [6]),
	.F(\top/processor/sha_core/n203_3 )
);
defparam \top/processor/sha_core/n203_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n204_s0  (
	.I0(\top/processor/sha_core/g [7]),
	.I1(\top/processor/sha_core/f [7]),
	.I2(\top/processor/sha_core/e [7]),
	.F(\top/processor/sha_core/n204_3 )
);
defparam \top/processor/sha_core/n204_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n205_s0  (
	.I0(\top/processor/sha_core/g [8]),
	.I1(\top/processor/sha_core/f [8]),
	.I2(\top/processor/sha_core/e [8]),
	.F(\top/processor/sha_core/n205_3 )
);
defparam \top/processor/sha_core/n205_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n206_s0  (
	.I0(\top/processor/sha_core/g [9]),
	.I1(\top/processor/sha_core/f [9]),
	.I2(\top/processor/sha_core/e [9]),
	.F(\top/processor/sha_core/n206_3 )
);
defparam \top/processor/sha_core/n206_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n207_s0  (
	.I0(\top/processor/sha_core/g [10]),
	.I1(\top/processor/sha_core/f [10]),
	.I2(\top/processor/sha_core/e [10]),
	.F(\top/processor/sha_core/n207_3 )
);
defparam \top/processor/sha_core/n207_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n208_s0  (
	.I0(\top/processor/sha_core/g [11]),
	.I1(\top/processor/sha_core/f [11]),
	.I2(\top/processor/sha_core/e [11]),
	.F(\top/processor/sha_core/n208_3 )
);
defparam \top/processor/sha_core/n208_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n209_s0  (
	.I0(\top/processor/sha_core/g [12]),
	.I1(\top/processor/sha_core/f [12]),
	.I2(\top/processor/sha_core/e [12]),
	.F(\top/processor/sha_core/n209_3 )
);
defparam \top/processor/sha_core/n209_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n210_s0  (
	.I0(\top/processor/sha_core/g [13]),
	.I1(\top/processor/sha_core/f [13]),
	.I2(\top/processor/sha_core/e [13]),
	.F(\top/processor/sha_core/n210_3 )
);
defparam \top/processor/sha_core/n210_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n211_s0  (
	.I0(\top/processor/sha_core/g [14]),
	.I1(\top/processor/sha_core/f [14]),
	.I2(\top/processor/sha_core/e [14]),
	.F(\top/processor/sha_core/n211_3 )
);
defparam \top/processor/sha_core/n211_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n212_s0  (
	.I0(\top/processor/sha_core/g [15]),
	.I1(\top/processor/sha_core/f [15]),
	.I2(\top/processor/sha_core/e [15]),
	.F(\top/processor/sha_core/n212_3 )
);
defparam \top/processor/sha_core/n212_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n213_s0  (
	.I0(\top/processor/sha_core/g [16]),
	.I1(\top/processor/sha_core/f [16]),
	.I2(\top/processor/sha_core/e [16]),
	.F(\top/processor/sha_core/n213_3 )
);
defparam \top/processor/sha_core/n213_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n214_s0  (
	.I0(\top/processor/sha_core/g [17]),
	.I1(\top/processor/sha_core/f [17]),
	.I2(\top/processor/sha_core/e [17]),
	.F(\top/processor/sha_core/n214_3 )
);
defparam \top/processor/sha_core/n214_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n215_s0  (
	.I0(\top/processor/sha_core/g [18]),
	.I1(\top/processor/sha_core/f [18]),
	.I2(\top/processor/sha_core/e [18]),
	.F(\top/processor/sha_core/n215_3 )
);
defparam \top/processor/sha_core/n215_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n216_s0  (
	.I0(\top/processor/sha_core/g [19]),
	.I1(\top/processor/sha_core/f [19]),
	.I2(\top/processor/sha_core/e [19]),
	.F(\top/processor/sha_core/n216_3 )
);
defparam \top/processor/sha_core/n216_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n217_s0  (
	.I0(\top/processor/sha_core/g [20]),
	.I1(\top/processor/sha_core/f [20]),
	.I2(\top/processor/sha_core/e [20]),
	.F(\top/processor/sha_core/n217_3 )
);
defparam \top/processor/sha_core/n217_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n218_s0  (
	.I0(\top/processor/sha_core/g [21]),
	.I1(\top/processor/sha_core/f [21]),
	.I2(\top/processor/sha_core/e [21]),
	.F(\top/processor/sha_core/n218_3 )
);
defparam \top/processor/sha_core/n218_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n219_s0  (
	.I0(\top/processor/sha_core/g [22]),
	.I1(\top/processor/sha_core/f [22]),
	.I2(\top/processor/sha_core/e [22]),
	.F(\top/processor/sha_core/n219_3 )
);
defparam \top/processor/sha_core/n219_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n220_s0  (
	.I0(\top/processor/sha_core/g [23]),
	.I1(\top/processor/sha_core/f [23]),
	.I2(\top/processor/sha_core/e [23]),
	.F(\top/processor/sha_core/n220_3 )
);
defparam \top/processor/sha_core/n220_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n221_s0  (
	.I0(\top/processor/sha_core/g [24]),
	.I1(\top/processor/sha_core/f [24]),
	.I2(\top/processor/sha_core/e [24]),
	.F(\top/processor/sha_core/n221_3 )
);
defparam \top/processor/sha_core/n221_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n222_s0  (
	.I0(\top/processor/sha_core/g [25]),
	.I1(\top/processor/sha_core/f [25]),
	.I2(\top/processor/sha_core/e [25]),
	.F(\top/processor/sha_core/n222_3 )
);
defparam \top/processor/sha_core/n222_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n223_s0  (
	.I0(\top/processor/sha_core/g [26]),
	.I1(\top/processor/sha_core/f [26]),
	.I2(\top/processor/sha_core/e [26]),
	.F(\top/processor/sha_core/n223_3 )
);
defparam \top/processor/sha_core/n223_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n224_s0  (
	.I0(\top/processor/sha_core/g [27]),
	.I1(\top/processor/sha_core/f [27]),
	.I2(\top/processor/sha_core/e [27]),
	.F(\top/processor/sha_core/n224_3 )
);
defparam \top/processor/sha_core/n224_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n225_s0  (
	.I0(\top/processor/sha_core/g [28]),
	.I1(\top/processor/sha_core/f [28]),
	.I2(\top/processor/sha_core/e [28]),
	.F(\top/processor/sha_core/n225_3 )
);
defparam \top/processor/sha_core/n225_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n226_s0  (
	.I0(\top/processor/sha_core/g [29]),
	.I1(\top/processor/sha_core/f [29]),
	.I2(\top/processor/sha_core/e [29]),
	.F(\top/processor/sha_core/n226_3 )
);
defparam \top/processor/sha_core/n226_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n227_s0  (
	.I0(\top/processor/sha_core/g [30]),
	.I1(\top/processor/sha_core/f [30]),
	.I2(\top/processor/sha_core/e [30]),
	.F(\top/processor/sha_core/n227_3 )
);
defparam \top/processor/sha_core/n227_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n228_s0  (
	.I0(\top/processor/sha_core/g [31]),
	.I1(\top/processor/sha_core/f [31]),
	.I2(\top/processor/sha_core/e [31]),
	.F(\top/processor/sha_core/n228_3 )
);
defparam \top/processor/sha_core/n228_s0 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n424_s0  (
	.I0(\top/processor/sha_core/a [2]),
	.I1(\top/processor/sha_core/a [13]),
	.I2(\top/processor/sha_core/a [22]),
	.F(\top/processor/sha_core/n424_3 )
);
defparam \top/processor/sha_core/n424_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n425_s0  (
	.I0(\top/processor/sha_core/a [3]),
	.I1(\top/processor/sha_core/a [14]),
	.I2(\top/processor/sha_core/a [23]),
	.F(\top/processor/sha_core/n425_3 )
);
defparam \top/processor/sha_core/n425_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n426_s0  (
	.I0(\top/processor/sha_core/a [4]),
	.I1(\top/processor/sha_core/a [15]),
	.I2(\top/processor/sha_core/a [24]),
	.F(\top/processor/sha_core/n426_3 )
);
defparam \top/processor/sha_core/n426_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n427_s0  (
	.I0(\top/processor/sha_core/a [5]),
	.I1(\top/processor/sha_core/a [16]),
	.I2(\top/processor/sha_core/a [25]),
	.F(\top/processor/sha_core/n427_3 )
);
defparam \top/processor/sha_core/n427_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n428_s0  (
	.I0(\top/processor/sha_core/a [6]),
	.I1(\top/processor/sha_core/a [17]),
	.I2(\top/processor/sha_core/a [26]),
	.F(\top/processor/sha_core/n428_3 )
);
defparam \top/processor/sha_core/n428_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n429_s0  (
	.I0(\top/processor/sha_core/a [7]),
	.I1(\top/processor/sha_core/a [18]),
	.I2(\top/processor/sha_core/a [27]),
	.F(\top/processor/sha_core/n429_3 )
);
defparam \top/processor/sha_core/n429_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n430_s0  (
	.I0(\top/processor/sha_core/a [8]),
	.I1(\top/processor/sha_core/a [19]),
	.I2(\top/processor/sha_core/a [28]),
	.F(\top/processor/sha_core/n430_3 )
);
defparam \top/processor/sha_core/n430_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n431_s0  (
	.I0(\top/processor/sha_core/a [9]),
	.I1(\top/processor/sha_core/a [20]),
	.I2(\top/processor/sha_core/a [29]),
	.F(\top/processor/sha_core/n431_3 )
);
defparam \top/processor/sha_core/n431_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n432_s0  (
	.I0(\top/processor/sha_core/a [10]),
	.I1(\top/processor/sha_core/a [21]),
	.I2(\top/processor/sha_core/a [30]),
	.F(\top/processor/sha_core/n432_3 )
);
defparam \top/processor/sha_core/n432_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n433_s0  (
	.I0(\top/processor/sha_core/a [11]),
	.I1(\top/processor/sha_core/a [22]),
	.I2(\top/processor/sha_core/a [31]),
	.F(\top/processor/sha_core/n433_3 )
);
defparam \top/processor/sha_core/n433_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n434_s0  (
	.I0(\top/processor/sha_core/a [12]),
	.I1(\top/processor/sha_core/a [23]),
	.I2(\top/processor/sha_core/a [0]),
	.F(\top/processor/sha_core/n434_3 )
);
defparam \top/processor/sha_core/n434_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n435_s0  (
	.I0(\top/processor/sha_core/a [13]),
	.I1(\top/processor/sha_core/a [24]),
	.I2(\top/processor/sha_core/a [1]),
	.F(\top/processor/sha_core/n435_3 )
);
defparam \top/processor/sha_core/n435_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n436_s0  (
	.I0(\top/processor/sha_core/a [2]),
	.I1(\top/processor/sha_core/a [14]),
	.I2(\top/processor/sha_core/a [25]),
	.F(\top/processor/sha_core/n436_3 )
);
defparam \top/processor/sha_core/n436_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n437_s0  (
	.I0(\top/processor/sha_core/a [3]),
	.I1(\top/processor/sha_core/a [15]),
	.I2(\top/processor/sha_core/a [26]),
	.F(\top/processor/sha_core/n437_3 )
);
defparam \top/processor/sha_core/n437_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n438_s0  (
	.I0(\top/processor/sha_core/a [4]),
	.I1(\top/processor/sha_core/a [16]),
	.I2(\top/processor/sha_core/a [27]),
	.F(\top/processor/sha_core/n438_3 )
);
defparam \top/processor/sha_core/n438_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n439_s0  (
	.I0(\top/processor/sha_core/a [5]),
	.I1(\top/processor/sha_core/a [17]),
	.I2(\top/processor/sha_core/a [28]),
	.F(\top/processor/sha_core/n439_3 )
);
defparam \top/processor/sha_core/n439_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n440_s0  (
	.I0(\top/processor/sha_core/a [6]),
	.I1(\top/processor/sha_core/a [18]),
	.I2(\top/processor/sha_core/a [29]),
	.F(\top/processor/sha_core/n440_3 )
);
defparam \top/processor/sha_core/n440_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n441_s0  (
	.I0(\top/processor/sha_core/a [7]),
	.I1(\top/processor/sha_core/a [19]),
	.I2(\top/processor/sha_core/a [30]),
	.F(\top/processor/sha_core/n441_3 )
);
defparam \top/processor/sha_core/n441_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n442_s0  (
	.I0(\top/processor/sha_core/a [8]),
	.I1(\top/processor/sha_core/a [20]),
	.I2(\top/processor/sha_core/a [31]),
	.F(\top/processor/sha_core/n442_3 )
);
defparam \top/processor/sha_core/n442_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n443_s0  (
	.I0(\top/processor/sha_core/a [9]),
	.I1(\top/processor/sha_core/a [21]),
	.I2(\top/processor/sha_core/a [0]),
	.F(\top/processor/sha_core/n443_3 )
);
defparam \top/processor/sha_core/n443_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n444_s0  (
	.I0(\top/processor/sha_core/a [10]),
	.I1(\top/processor/sha_core/a [22]),
	.I2(\top/processor/sha_core/a [1]),
	.F(\top/processor/sha_core/n444_3 )
);
defparam \top/processor/sha_core/n444_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n445_s0  (
	.I0(\top/processor/sha_core/a [2]),
	.I1(\top/processor/sha_core/a [11]),
	.I2(\top/processor/sha_core/a [23]),
	.F(\top/processor/sha_core/n445_3 )
);
defparam \top/processor/sha_core/n445_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n446_s0  (
	.I0(\top/processor/sha_core/a [3]),
	.I1(\top/processor/sha_core/a [12]),
	.I2(\top/processor/sha_core/a [24]),
	.F(\top/processor/sha_core/n446_3 )
);
defparam \top/processor/sha_core/n446_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n447_s0  (
	.I0(\top/processor/sha_core/a [13]),
	.I1(\top/processor/sha_core/a [4]),
	.I2(\top/processor/sha_core/a [25]),
	.F(\top/processor/sha_core/n447_3 )
);
defparam \top/processor/sha_core/n447_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n448_s0  (
	.I0(\top/processor/sha_core/a [14]),
	.I1(\top/processor/sha_core/a [5]),
	.I2(\top/processor/sha_core/a [26]),
	.F(\top/processor/sha_core/n448_3 )
);
defparam \top/processor/sha_core/n448_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n449_s0  (
	.I0(\top/processor/sha_core/a [15]),
	.I1(\top/processor/sha_core/a [6]),
	.I2(\top/processor/sha_core/a [27]),
	.F(\top/processor/sha_core/n449_3 )
);
defparam \top/processor/sha_core/n449_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n450_s0  (
	.I0(\top/processor/sha_core/a [16]),
	.I1(\top/processor/sha_core/a [7]),
	.I2(\top/processor/sha_core/a [28]),
	.F(\top/processor/sha_core/n450_3 )
);
defparam \top/processor/sha_core/n450_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n451_s0  (
	.I0(\top/processor/sha_core/a [17]),
	.I1(\top/processor/sha_core/a [8]),
	.I2(\top/processor/sha_core/a [29]),
	.F(\top/processor/sha_core/n451_3 )
);
defparam \top/processor/sha_core/n451_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n452_s0  (
	.I0(\top/processor/sha_core/a [18]),
	.I1(\top/processor/sha_core/a [9]),
	.I2(\top/processor/sha_core/a [30]),
	.F(\top/processor/sha_core/n452_3 )
);
defparam \top/processor/sha_core/n452_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n453_s0  (
	.I0(\top/processor/sha_core/a [19]),
	.I1(\top/processor/sha_core/a [10]),
	.I2(\top/processor/sha_core/a [31]),
	.F(\top/processor/sha_core/n453_3 )
);
defparam \top/processor/sha_core/n453_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n454_s0  (
	.I0(\top/processor/sha_core/a [20]),
	.I1(\top/processor/sha_core/a [11]),
	.I2(\top/processor/sha_core/a [0]),
	.F(\top/processor/sha_core/n454_3 )
);
defparam \top/processor/sha_core/n454_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n455_s0  (
	.I0(\top/processor/sha_core/a [21]),
	.I1(\top/processor/sha_core/a [12]),
	.I2(\top/processor/sha_core/a [1]),
	.F(\top/processor/sha_core/n455_3 )
);
defparam \top/processor/sha_core/n455_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n584_s0  (
	.I0(\top/processor/sha_core/a [0]),
	.I1(\top/processor/sha_core/b [0]),
	.I2(\top/processor/sha_core/c [0]),
	.F(\top/processor/sha_core/n584_3 )
);
defparam \top/processor/sha_core/n584_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n585_s0  (
	.I0(\top/processor/sha_core/a [1]),
	.I1(\top/processor/sha_core/b [1]),
	.I2(\top/processor/sha_core/c [1]),
	.F(\top/processor/sha_core/n585_3 )
);
defparam \top/processor/sha_core/n585_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n586_s0  (
	.I0(\top/processor/sha_core/a [2]),
	.I1(\top/processor/sha_core/b [2]),
	.I2(\top/processor/sha_core/c [2]),
	.F(\top/processor/sha_core/n586_3 )
);
defparam \top/processor/sha_core/n586_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n587_s0  (
	.I0(\top/processor/sha_core/a [3]),
	.I1(\top/processor/sha_core/b [3]),
	.I2(\top/processor/sha_core/c [3]),
	.F(\top/processor/sha_core/n587_3 )
);
defparam \top/processor/sha_core/n587_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n588_s0  (
	.I0(\top/processor/sha_core/a [4]),
	.I1(\top/processor/sha_core/b [4]),
	.I2(\top/processor/sha_core/c [4]),
	.F(\top/processor/sha_core/n588_3 )
);
defparam \top/processor/sha_core/n588_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n589_s0  (
	.I0(\top/processor/sha_core/a [5]),
	.I1(\top/processor/sha_core/b [5]),
	.I2(\top/processor/sha_core/c [5]),
	.F(\top/processor/sha_core/n589_3 )
);
defparam \top/processor/sha_core/n589_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n590_s0  (
	.I0(\top/processor/sha_core/a [6]),
	.I1(\top/processor/sha_core/b [6]),
	.I2(\top/processor/sha_core/c [6]),
	.F(\top/processor/sha_core/n590_3 )
);
defparam \top/processor/sha_core/n590_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n591_s0  (
	.I0(\top/processor/sha_core/a [7]),
	.I1(\top/processor/sha_core/b [7]),
	.I2(\top/processor/sha_core/c [7]),
	.F(\top/processor/sha_core/n591_3 )
);
defparam \top/processor/sha_core/n591_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n592_s0  (
	.I0(\top/processor/sha_core/a [8]),
	.I1(\top/processor/sha_core/b [8]),
	.I2(\top/processor/sha_core/c [8]),
	.F(\top/processor/sha_core/n592_3 )
);
defparam \top/processor/sha_core/n592_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n593_s0  (
	.I0(\top/processor/sha_core/a [9]),
	.I1(\top/processor/sha_core/b [9]),
	.I2(\top/processor/sha_core/c [9]),
	.F(\top/processor/sha_core/n593_3 )
);
defparam \top/processor/sha_core/n593_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n594_s0  (
	.I0(\top/processor/sha_core/a [10]),
	.I1(\top/processor/sha_core/b [10]),
	.I2(\top/processor/sha_core/c [10]),
	.F(\top/processor/sha_core/n594_3 )
);
defparam \top/processor/sha_core/n594_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n595_s0  (
	.I0(\top/processor/sha_core/a [11]),
	.I1(\top/processor/sha_core/b [11]),
	.I2(\top/processor/sha_core/c [11]),
	.F(\top/processor/sha_core/n595_3 )
);
defparam \top/processor/sha_core/n595_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n596_s0  (
	.I0(\top/processor/sha_core/a [12]),
	.I1(\top/processor/sha_core/b [12]),
	.I2(\top/processor/sha_core/c [12]),
	.F(\top/processor/sha_core/n596_3 )
);
defparam \top/processor/sha_core/n596_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n597_s0  (
	.I0(\top/processor/sha_core/a [13]),
	.I1(\top/processor/sha_core/b [13]),
	.I2(\top/processor/sha_core/c [13]),
	.F(\top/processor/sha_core/n597_3 )
);
defparam \top/processor/sha_core/n597_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n598_s0  (
	.I0(\top/processor/sha_core/a [14]),
	.I1(\top/processor/sha_core/b [14]),
	.I2(\top/processor/sha_core/c [14]),
	.F(\top/processor/sha_core/n598_3 )
);
defparam \top/processor/sha_core/n598_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n599_s0  (
	.I0(\top/processor/sha_core/a [15]),
	.I1(\top/processor/sha_core/b [15]),
	.I2(\top/processor/sha_core/c [15]),
	.F(\top/processor/sha_core/n599_3 )
);
defparam \top/processor/sha_core/n599_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n600_s0  (
	.I0(\top/processor/sha_core/a [16]),
	.I1(\top/processor/sha_core/b [16]),
	.I2(\top/processor/sha_core/c [16]),
	.F(\top/processor/sha_core/n600_3 )
);
defparam \top/processor/sha_core/n600_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n601_s0  (
	.I0(\top/processor/sha_core/a [17]),
	.I1(\top/processor/sha_core/b [17]),
	.I2(\top/processor/sha_core/c [17]),
	.F(\top/processor/sha_core/n601_3 )
);
defparam \top/processor/sha_core/n601_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n602_s0  (
	.I0(\top/processor/sha_core/a [18]),
	.I1(\top/processor/sha_core/b [18]),
	.I2(\top/processor/sha_core/c [18]),
	.F(\top/processor/sha_core/n602_3 )
);
defparam \top/processor/sha_core/n602_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n603_s0  (
	.I0(\top/processor/sha_core/a [19]),
	.I1(\top/processor/sha_core/b [19]),
	.I2(\top/processor/sha_core/c [19]),
	.F(\top/processor/sha_core/n603_3 )
);
defparam \top/processor/sha_core/n603_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n604_s0  (
	.I0(\top/processor/sha_core/a [20]),
	.I1(\top/processor/sha_core/b [20]),
	.I2(\top/processor/sha_core/c [20]),
	.F(\top/processor/sha_core/n604_3 )
);
defparam \top/processor/sha_core/n604_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n605_s0  (
	.I0(\top/processor/sha_core/a [21]),
	.I1(\top/processor/sha_core/b [21]),
	.I2(\top/processor/sha_core/c [21]),
	.F(\top/processor/sha_core/n605_3 )
);
defparam \top/processor/sha_core/n605_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n606_s0  (
	.I0(\top/processor/sha_core/a [22]),
	.I1(\top/processor/sha_core/b [22]),
	.I2(\top/processor/sha_core/c [22]),
	.F(\top/processor/sha_core/n606_3 )
);
defparam \top/processor/sha_core/n606_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n607_s0  (
	.I0(\top/processor/sha_core/a [23]),
	.I1(\top/processor/sha_core/b [23]),
	.I2(\top/processor/sha_core/c [23]),
	.F(\top/processor/sha_core/n607_3 )
);
defparam \top/processor/sha_core/n607_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n608_s0  (
	.I0(\top/processor/sha_core/a [24]),
	.I1(\top/processor/sha_core/b [24]),
	.I2(\top/processor/sha_core/c [24]),
	.F(\top/processor/sha_core/n608_3 )
);
defparam \top/processor/sha_core/n608_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n609_s0  (
	.I0(\top/processor/sha_core/a [25]),
	.I1(\top/processor/sha_core/b [25]),
	.I2(\top/processor/sha_core/c [25]),
	.F(\top/processor/sha_core/n609_3 )
);
defparam \top/processor/sha_core/n609_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n610_s0  (
	.I0(\top/processor/sha_core/a [26]),
	.I1(\top/processor/sha_core/b [26]),
	.I2(\top/processor/sha_core/c [26]),
	.F(\top/processor/sha_core/n610_3 )
);
defparam \top/processor/sha_core/n610_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n611_s0  (
	.I0(\top/processor/sha_core/a [27]),
	.I1(\top/processor/sha_core/b [27]),
	.I2(\top/processor/sha_core/c [27]),
	.F(\top/processor/sha_core/n611_3 )
);
defparam \top/processor/sha_core/n611_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n612_s0  (
	.I0(\top/processor/sha_core/a [28]),
	.I1(\top/processor/sha_core/b [28]),
	.I2(\top/processor/sha_core/c [28]),
	.F(\top/processor/sha_core/n612_3 )
);
defparam \top/processor/sha_core/n612_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n613_s0  (
	.I0(\top/processor/sha_core/a [29]),
	.I1(\top/processor/sha_core/b [29]),
	.I2(\top/processor/sha_core/c [29]),
	.F(\top/processor/sha_core/n613_3 )
);
defparam \top/processor/sha_core/n613_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n614_s0  (
	.I0(\top/processor/sha_core/a [30]),
	.I1(\top/processor/sha_core/b [30]),
	.I2(\top/processor/sha_core/c [30]),
	.F(\top/processor/sha_core/n614_3 )
);
defparam \top/processor/sha_core/n614_s0 .INIT=8'hE8;
LUT3 \top/processor/sha_core/n615_s0  (
	.I0(\top/processor/sha_core/a [31]),
	.I1(\top/processor/sha_core/b [31]),
	.I2(\top/processor/sha_core/c [31]),
	.F(\top/processor/sha_core/n615_3 )
);
defparam \top/processor/sha_core/n615_s0 .INIT=8'hE8;
LUT2 \top/processor/sha_core/n3543_s0  (
	.I0(\top/processor/sha_core/n3511_193 ),
	.I1(\top/processor/sha_core/n3509_193 ),
	.F(\top/processor/sha_core/n3543_3 )
);
defparam \top/processor/sha_core/n3543_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3545_s0  (
	.I0(\top/processor/sha_core/n3509_193 ),
	.I1(\top/processor/sha_core/n3507_193 ),
	.F(\top/processor/sha_core/n3545_3 )
);
defparam \top/processor/sha_core/n3545_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3546_s0  (
	.I0(\top/processor/sha_core/n3508_193 ),
	.I1(\top/processor/sha_core/n3506_193 ),
	.F(\top/processor/sha_core/n3546_3 )
);
defparam \top/processor/sha_core/n3546_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3547_s0  (
	.I0(\top/processor/sha_core/n3507_193 ),
	.I1(\top/processor/sha_core/n3505_193 ),
	.F(\top/processor/sha_core/n3547_3 )
);
defparam \top/processor/sha_core/n3547_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3548_s0  (
	.I0(\top/processor/sha_core/n3506_193 ),
	.I1(\top/processor/sha_core/n3504_193 ),
	.F(\top/processor/sha_core/n3548_3 )
);
defparam \top/processor/sha_core/n3548_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3549_s0  (
	.I0(\top/processor/sha_core/n3505_193 ),
	.I1(\top/processor/sha_core/n3503_193 ),
	.F(\top/processor/sha_core/n3549_3 )
);
defparam \top/processor/sha_core/n3549_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3550_s0  (
	.I0(\top/processor/sha_core/n3502_193 ),
	.I1(\top/processor/sha_core/n3504_193 ),
	.F(\top/processor/sha_core/n3550_3 )
);
defparam \top/processor/sha_core/n3550_s0 .INIT=4'h6;
LUT2 \top/processor/sha_core/n3551_s0  (
	.I0(\top/processor/sha_core/n3501_193 ),
	.I1(\top/processor/sha_core/n3503_193 ),
	.F(\top/processor/sha_core/n3551_3 )
);
defparam \top/processor/sha_core/n3551_s0 .INIT=4'h6;
LUT3 \top/processor/sha_core/n3552_s0  (
	.I0(\top/processor/sha_core/n3502_193 ),
	.I1(\top/processor/sha_core/n3500_193 ),
	.I2(\top/processor/sha_core/n3509_193 ),
	.F(\top/processor/sha_core/n3552_3 )
);
defparam \top/processor/sha_core/n3552_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3553_s0  (
	.I0(\top/processor/sha_core/n3501_193 ),
	.I1(\top/processor/sha_core/n3499_193 ),
	.I2(\top/processor/sha_core/n3508_193 ),
	.F(\top/processor/sha_core/n3553_3 )
);
defparam \top/processor/sha_core/n3553_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3554_s0  (
	.I0(\top/processor/sha_core/n3500_193 ),
	.I1(\top/processor/sha_core/n3498_193 ),
	.I2(\top/processor/sha_core/n3507_193 ),
	.F(\top/processor/sha_core/n3554_3 )
);
defparam \top/processor/sha_core/n3554_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3555_s0  (
	.I0(\top/processor/sha_core/n3499_193 ),
	.I1(\top/processor/sha_core/n3497_193 ),
	.I2(\top/processor/sha_core/n3506_193 ),
	.F(\top/processor/sha_core/n3555_3 )
);
defparam \top/processor/sha_core/n3555_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3556_s0  (
	.I0(\top/processor/sha_core/n3498_193 ),
	.I1(\top/processor/sha_core/n3496_193 ),
	.I2(\top/processor/sha_core/n3505_193 ),
	.F(\top/processor/sha_core/n3556_3 )
);
defparam \top/processor/sha_core/n3556_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3557_s0  (
	.I0(\top/processor/sha_core/n3497_193 ),
	.I1(\top/processor/sha_core/n3495_193 ),
	.I2(\top/processor/sha_core/n3504_193 ),
	.F(\top/processor/sha_core/n3557_3 )
);
defparam \top/processor/sha_core/n3557_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3558_s0  (
	.I0(\top/processor/sha_core/n3496_193 ),
	.I1(\top/processor/sha_core/n3494_194 ),
	.I2(\top/processor/sha_core/n3503_193 ),
	.F(\top/processor/sha_core/n3558_3 )
);
defparam \top/processor/sha_core/n3558_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3559_s0  (
	.I0(\top/processor/sha_core/n3502_193 ),
	.I1(\top/processor/sha_core/n3495_193 ),
	.I2(\top/processor/sha_core/n3493_193 ),
	.F(\top/processor/sha_core/n3559_3 )
);
defparam \top/processor/sha_core/n3559_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3560_s0  (
	.I0(\top/processor/sha_core/n3501_193 ),
	.I1(\top/processor/sha_core/n3494_194 ),
	.I2(\top/processor/sha_core/n3492_193 ),
	.F(\top/processor/sha_core/n3560_3 )
);
defparam \top/processor/sha_core/n3560_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3561_s0  (
	.I0(\top/processor/sha_core/n3500_193 ),
	.I1(\top/processor/sha_core/n3493_193 ),
	.I2(\top/processor/sha_core/n3491_193 ),
	.F(\top/processor/sha_core/n3561_3 )
);
defparam \top/processor/sha_core/n3561_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3562_s0  (
	.I0(\top/processor/sha_core/n3499_193 ),
	.I1(\top/processor/sha_core/n3492_193 ),
	.I2(\top/processor/sha_core/n3490_193 ),
	.F(\top/processor/sha_core/n3562_3 )
);
defparam \top/processor/sha_core/n3562_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3563_s0  (
	.I0(\top/processor/sha_core/n3498_193 ),
	.I1(\top/processor/sha_core/n3491_193 ),
	.I2(\top/processor/sha_core/n3489_193 ),
	.F(\top/processor/sha_core/n3563_3 )
);
defparam \top/processor/sha_core/n3563_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3564_s0  (
	.I0(\top/processor/sha_core/n3497_193 ),
	.I1(\top/processor/sha_core/n3490_193 ),
	.I2(\top/processor/sha_core/n3488_193 ),
	.F(\top/processor/sha_core/n3564_3 )
);
defparam \top/processor/sha_core/n3564_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3565_s0  (
	.I0(\top/processor/sha_core/n3496_193 ),
	.I1(\top/processor/sha_core/n3489_193 ),
	.I2(\top/processor/sha_core/n3519_193 ),
	.F(\top/processor/sha_core/n3565_3 )
);
defparam \top/processor/sha_core/n3565_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3566_s0  (
	.I0(\top/processor/sha_core/n3495_193 ),
	.I1(\top/processor/sha_core/n3488_193 ),
	.I2(\top/processor/sha_core/n3518_193 ),
	.F(\top/processor/sha_core/n3566_3 )
);
defparam \top/processor/sha_core/n3566_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3567_s0  (
	.I0(\top/processor/sha_core/n3494_194 ),
	.I1(\top/processor/sha_core/n3519_193 ),
	.I2(\top/processor/sha_core/n3517_193 ),
	.F(\top/processor/sha_core/n3567_3 )
);
defparam \top/processor/sha_core/n3567_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3568_s0  (
	.I0(\top/processor/sha_core/n3493_193 ),
	.I1(\top/processor/sha_core/n3518_193 ),
	.I2(\top/processor/sha_core/n3516_193 ),
	.F(\top/processor/sha_core/n3568_3 )
);
defparam \top/processor/sha_core/n3568_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3569_s0  (
	.I0(\top/processor/sha_core/n3492_193 ),
	.I1(\top/processor/sha_core/n3517_193 ),
	.I2(\top/processor/sha_core/n3515_193 ),
	.F(\top/processor/sha_core/n3569_3 )
);
defparam \top/processor/sha_core/n3569_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3570_s0  (
	.I0(\top/processor/sha_core/n3491_193 ),
	.I1(\top/processor/sha_core/n3516_193 ),
	.I2(\top/processor/sha_core/n3514_193 ),
	.F(\top/processor/sha_core/n3570_3 )
);
defparam \top/processor/sha_core/n3570_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3571_s0  (
	.I0(\top/processor/sha_core/n3490_193 ),
	.I1(\top/processor/sha_core/n3515_193 ),
	.I2(\top/processor/sha_core/n3513_193 ),
	.F(\top/processor/sha_core/n3571_3 )
);
defparam \top/processor/sha_core/n3571_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3572_s0  (
	.I0(\top/processor/sha_core/n3489_193 ),
	.I1(\top/processor/sha_core/n3514_193 ),
	.I2(\top/processor/sha_core/n3512_193 ),
	.F(\top/processor/sha_core/n3572_3 )
);
defparam \top/processor/sha_core/n3572_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3573_s0  (
	.I0(\top/processor/sha_core/n3488_193 ),
	.I1(\top/processor/sha_core/n3513_193 ),
	.I2(\top/processor/sha_core/n3511_193 ),
	.F(\top/processor/sha_core/n3573_3 )
);
defparam \top/processor/sha_core/n3573_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3769_s0  (
	.I0(\top/processor/sha_core/n3769_4 ),
	.I1(\top/processor/sha_core/n3769_5 ),
	.I2(\top/processor/sha_core/n3769_6 ),
	.F(\top/processor/sha_core/n3769_3 )
);
defparam \top/processor/sha_core/n3769_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3770_s0  (
	.I0(\top/processor/sha_core/n3766_5 ),
	.I1(\top/processor/sha_core/n3770_4 ),
	.I2(\top/processor/sha_core/n3770_5 ),
	.F(\top/processor/sha_core/n3770_3 )
);
defparam \top/processor/sha_core/n3770_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3771_s0  (
	.I0(\top/processor/sha_core/n3767_5 ),
	.I1(\top/processor/sha_core/n3771_4 ),
	.I2(\top/processor/sha_core/n3771_5 ),
	.F(\top/processor/sha_core/n3771_3 )
);
defparam \top/processor/sha_core/n3771_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3772_s0  (
	.I0(\top/processor/sha_core/n3768_5 ),
	.I1(\top/processor/sha_core/n3772_4 ),
	.I2(\top/processor/sha_core/n3772_5 ),
	.F(\top/processor/sha_core/n3772_3 )
);
defparam \top/processor/sha_core/n3772_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3773_s0  (
	.I0(\top/processor/sha_core/n3769_5 ),
	.I1(\top/processor/sha_core/n3773_4 ),
	.I2(\top/processor/sha_core/n3773_5 ),
	.F(\top/processor/sha_core/n3773_3 )
);
defparam \top/processor/sha_core/n3773_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3774_s0  (
	.I0(\top/processor/sha_core/n3770_5 ),
	.I1(\top/processor/sha_core/n3774_4 ),
	.I2(\top/processor/sha_core/n3774_5 ),
	.F(\top/processor/sha_core/n3774_3 )
);
defparam \top/processor/sha_core/n3774_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3775_s0  (
	.I0(\top/processor/sha_core/n3771_5 ),
	.I1(\top/processor/sha_core/n3775_4 ),
	.I2(\top/processor/sha_core/n3775_5 ),
	.F(\top/processor/sha_core/n3775_3 )
);
defparam \top/processor/sha_core/n3775_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3776_s0  (
	.I0(\top/processor/sha_core/n3772_4 ),
	.I1(\top/processor/sha_core/n3776_4 ),
	.I2(\top/processor/sha_core/n3776_5 ),
	.F(\top/processor/sha_core/n3776_3 )
);
defparam \top/processor/sha_core/n3776_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3777_s0  (
	.I0(\top/processor/sha_core/n3766_4 ),
	.I1(\top/processor/sha_core/n3773_4 ),
	.I2(\top/processor/sha_core/n3777_4 ),
	.F(\top/processor/sha_core/n3777_3 )
);
defparam \top/processor/sha_core/n3777_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3778_s0  (
	.I0(\top/processor/sha_core/n3767_4 ),
	.I1(\top/processor/sha_core/n3774_4 ),
	.I2(\top/processor/sha_core/n3778_4 ),
	.F(\top/processor/sha_core/n3778_3 )
);
defparam \top/processor/sha_core/n3778_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3779_s0  (
	.I0(\top/processor/sha_core/n3768_4 ),
	.I1(\top/processor/sha_core/n3775_4 ),
	.I2(\top/processor/sha_core/n3779_4 ),
	.F(\top/processor/sha_core/n3779_3 )
);
defparam \top/processor/sha_core/n3779_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3780_s0  (
	.I0(\top/processor/sha_core/n3769_4 ),
	.I1(\top/processor/sha_core/n3776_5 ),
	.I2(\top/processor/sha_core/n3780_4 ),
	.F(\top/processor/sha_core/n3780_3 )
);
defparam \top/processor/sha_core/n3780_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3781_s0  (
	.I0(\top/processor/sha_core/n3766_4 ),
	.I1(\top/processor/sha_core/n3770_4 ),
	.I2(\top/processor/sha_core/n3781_4 ),
	.F(\top/processor/sha_core/n3781_3 )
);
defparam \top/processor/sha_core/n3781_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3782_s0  (
	.I0(\top/processor/sha_core/n3767_4 ),
	.I1(\top/processor/sha_core/n3771_4 ),
	.I2(\top/processor/sha_core/n3782_4 ),
	.F(\top/processor/sha_core/n3782_3 )
);
defparam \top/processor/sha_core/n3782_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3783_s0  (
	.I0(\top/processor/sha_core/n3768_4 ),
	.I1(\top/processor/sha_core/n3772_5 ),
	.I2(\top/processor/sha_core/n3783_4 ),
	.F(\top/processor/sha_core/n3783_3 )
);
defparam \top/processor/sha_core/n3783_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3784_s0  (
	.I0(\top/processor/sha_core/n3769_4 ),
	.I1(\top/processor/sha_core/n3773_5 ),
	.I2(\top/processor/sha_core/n3784_4 ),
	.F(\top/processor/sha_core/n3784_3 )
);
defparam \top/processor/sha_core/n3784_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3785_s0  (
	.I0(\top/processor/sha_core/n3770_4 ),
	.I1(\top/processor/sha_core/n3774_5 ),
	.I2(\top/processor/sha_core/n3785_4 ),
	.F(\top/processor/sha_core/n3785_3 )
);
defparam \top/processor/sha_core/n3785_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3786_s0  (
	.I0(\top/processor/sha_core/n3769_6 ),
	.I1(\top/processor/sha_core/n3771_4 ),
	.I2(\top/processor/sha_core/n3775_5 ),
	.F(\top/processor/sha_core/n3786_3 )
);
defparam \top/processor/sha_core/n3786_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3787_s0  (
	.I0(\top/processor/sha_core/n3766_5 ),
	.I1(\top/processor/sha_core/n3772_5 ),
	.I2(\top/processor/sha_core/n3776_4 ),
	.F(\top/processor/sha_core/n3787_3 )
);
defparam \top/processor/sha_core/n3787_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3788_s0  (
	.I0(\top/processor/sha_core/n3767_5 ),
	.I1(\top/processor/sha_core/n3773_5 ),
	.I2(\top/processor/sha_core/n3777_4 ),
	.F(\top/processor/sha_core/n3788_3 )
);
defparam \top/processor/sha_core/n3788_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3789_s0  (
	.I0(\top/processor/sha_core/n3768_5 ),
	.I1(\top/processor/sha_core/n3774_5 ),
	.I2(\top/processor/sha_core/n3778_4 ),
	.F(\top/processor/sha_core/n3789_3 )
);
defparam \top/processor/sha_core/n3789_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3790_s0  (
	.I0(\top/processor/sha_core/n3769_5 ),
	.I1(\top/processor/sha_core/n3775_5 ),
	.I2(\top/processor/sha_core/n3779_4 ),
	.F(\top/processor/sha_core/n3790_3 )
);
defparam \top/processor/sha_core/n3790_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3791_s0  (
	.I0(\top/processor/sha_core/n3770_5 ),
	.I1(\top/processor/sha_core/n3776_4 ),
	.I2(\top/processor/sha_core/n3780_4 ),
	.F(\top/processor/sha_core/n3791_3 )
);
defparam \top/processor/sha_core/n3791_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3792_s0  (
	.I0(\top/processor/sha_core/n3771_5 ),
	.I1(\top/processor/sha_core/n3777_4 ),
	.I2(\top/processor/sha_core/n3781_4 ),
	.F(\top/processor/sha_core/n3792_3 )
);
defparam \top/processor/sha_core/n3792_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3793_s0  (
	.I0(\top/processor/sha_core/n3772_4 ),
	.I1(\top/processor/sha_core/n3778_4 ),
	.I2(\top/processor/sha_core/n3782_4 ),
	.F(\top/processor/sha_core/n3793_3 )
);
defparam \top/processor/sha_core/n3793_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3794_s0  (
	.I0(\top/processor/sha_core/n3773_4 ),
	.I1(\top/processor/sha_core/n3779_4 ),
	.I2(\top/processor/sha_core/n3783_4 ),
	.F(\top/processor/sha_core/n3794_3 )
);
defparam \top/processor/sha_core/n3794_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3795_s0  (
	.I0(\top/processor/sha_core/n3774_4 ),
	.I1(\top/processor/sha_core/n3780_4 ),
	.I2(\top/processor/sha_core/n3784_4 ),
	.F(\top/processor/sha_core/n3795_3 )
);
defparam \top/processor/sha_core/n3795_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3796_s0  (
	.I0(\top/processor/sha_core/n3775_4 ),
	.I1(\top/processor/sha_core/n3781_4 ),
	.I2(\top/processor/sha_core/n3785_4 ),
	.F(\top/processor/sha_core/n3796_3 )
);
defparam \top/processor/sha_core/n3796_s0 .INIT=8'h96;
LUT3 \top/processor/sha_core/n3797_s0  (
	.I0(\top/processor/sha_core/n3769_6 ),
	.I1(\top/processor/sha_core/n3776_5 ),
	.I2(\top/processor/sha_core/n3782_4 ),
	.F(\top/processor/sha_core/n3797_3 )
);
defparam \top/processor/sha_core/n3797_s0 .INIT=8'h96;
LUT4 \top/processor/sha_core/n8430_s0  (
	.I0(\top/processor/sha_core/n8430_4 ),
	.I1(\top/processor/sha_core/n8430_5 ),
	.I2(\top/processor/sha_core/n3893_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8430_3 )
);
defparam \top/processor/sha_core/n8430_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8431_s0  (
	.I0(\top/processor/sha_core/n8431_4 ),
	.I1(\top/processor/sha_core/n8431_5 ),
	.I2(\top/processor/sha_core/n3894_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8431_3 )
);
defparam \top/processor/sha_core/n8431_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8432_s0  (
	.I0(\top/processor/sha_core/n8432_4 ),
	.I1(\top/processor/sha_core/n8432_5 ),
	.I2(\top/processor/sha_core/n3895_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8432_3 )
);
defparam \top/processor/sha_core/n8432_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8433_s0  (
	.I0(\top/processor/sha_core/n8433_4 ),
	.I1(\top/processor/sha_core/n8433_5 ),
	.I2(\top/processor/sha_core/n3896_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8433_3 )
);
defparam \top/processor/sha_core/n8433_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8434_s0  (
	.I0(\top/processor/sha_core/n8434_4 ),
	.I1(\top/processor/sha_core/n8434_5 ),
	.I2(\top/processor/sha_core/n3897_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8434_3 )
);
defparam \top/processor/sha_core/n8434_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8435_s0  (
	.I0(\top/processor/sha_core/n8435_4 ),
	.I1(\top/processor/sha_core/n8435_5 ),
	.I2(\top/processor/sha_core/n3898_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8435_3 )
);
defparam \top/processor/sha_core/n8435_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8436_s0  (
	.I0(\top/processor/sha_core/n8436_4 ),
	.I1(\top/processor/sha_core/n8436_5 ),
	.I2(\top/processor/sha_core/n3899_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8436_3 )
);
defparam \top/processor/sha_core/n8436_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8437_s0  (
	.I0(\top/processor/sha_core/n8437_4 ),
	.I1(\top/processor/sha_core/n8437_5 ),
	.I2(\top/processor/sha_core/n3900_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8437_3 )
);
defparam \top/processor/sha_core/n8437_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8438_s0  (
	.I0(\top/processor/sha_core/n8438_4 ),
	.I1(\top/processor/sha_core/n8438_5 ),
	.I2(\top/processor/sha_core/n3901_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8438_3 )
);
defparam \top/processor/sha_core/n8438_s0 .INIT=16'h77F0;
LUT3 \top/processor/sha_core/n8439_s0  (
	.I0(\top/processor/sha_core/n3902_5 ),
	.I1(\top/processor/sha_core/n8439_4 ),
	.I2(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8439_3 )
);
defparam \top/processor/sha_core/n8439_s0 .INIT=8'h3A;
LUT4 \top/processor/sha_core/n8440_s0  (
	.I0(\top/processor/sha_core/n8440_4 ),
	.I1(\top/processor/sha_core/n8440_5 ),
	.I2(\top/processor/sha_core/n3903_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8440_3 )
);
defparam \top/processor/sha_core/n8440_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8441_s0  (
	.I0(\top/processor/sha_core/n8441_4 ),
	.I1(\top/processor/sha_core/n8441_5 ),
	.I2(\top/processor/sha_core/n3904_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8441_3 )
);
defparam \top/processor/sha_core/n8441_s0 .INIT=16'h77F0;
LUT3 \top/processor/sha_core/n8442_s0  (
	.I0(\top/processor/sha_core/n8442_4 ),
	.I1(\top/processor/sha_core/n3905_5 ),
	.I2(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8442_3 )
);
defparam \top/processor/sha_core/n8442_s0 .INIT=8'h5C;
LUT4 \top/processor/sha_core/n8443_s0  (
	.I0(\top/processor/sha_core/n8443_4 ),
	.I1(\top/processor/sha_core/n8443_5 ),
	.I2(\top/processor/sha_core/n3906_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8443_3 )
);
defparam \top/processor/sha_core/n8443_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8444_s0  (
	.I0(\top/processor/sha_core/n8444_4 ),
	.I1(\top/processor/sha_core/n8444_5 ),
	.I2(\top/processor/sha_core/n3907_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8444_3 )
);
defparam \top/processor/sha_core/n8444_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8445_s0  (
	.I0(\top/processor/sha_core/n8445_4 ),
	.I1(\top/processor/sha_core/n8445_5 ),
	.I2(\top/processor/sha_core/n3908_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8445_3 )
);
defparam \top/processor/sha_core/n8445_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8446_s0  (
	.I0(\top/processor/sha_core/n8446_4 ),
	.I1(\top/processor/sha_core/n8446_5 ),
	.I2(\top/processor/sha_core/n3909_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8446_3 )
);
defparam \top/processor/sha_core/n8446_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8447_s0  (
	.I0(\top/processor/sha_core/n8447_4 ),
	.I1(\top/processor/sha_core/n8447_5 ),
	.I2(\top/processor/sha_core/n3910_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8447_3 )
);
defparam \top/processor/sha_core/n8447_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8448_s0  (
	.I0(\top/processor/sha_core/n8448_4 ),
	.I1(\top/processor/sha_core/n8448_5 ),
	.I2(\top/processor/sha_core/n3911_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8448_3 )
);
defparam \top/processor/sha_core/n8448_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8449_s0  (
	.I0(\top/processor/sha_core/n8449_4 ),
	.I1(\top/processor/sha_core/n8449_5 ),
	.I2(\top/processor/sha_core/n3912_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8449_3 )
);
defparam \top/processor/sha_core/n8449_s0 .INIT=16'h77F0;
LUT3 \top/processor/sha_core/n8450_s0  (
	.I0(\top/processor/sha_core/n8450_4 ),
	.I1(\top/processor/sha_core/n3913_5 ),
	.I2(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8450_3 )
);
defparam \top/processor/sha_core/n8450_s0 .INIT=8'h5C;
LUT4 \top/processor/sha_core/n8451_s0  (
	.I0(\top/processor/sha_core/n8451_4 ),
	.I1(\top/processor/sha_core/n8451_5 ),
	.I2(\top/processor/sha_core/n3914_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8451_3 )
);
defparam \top/processor/sha_core/n8451_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8452_s0  (
	.I0(\top/processor/sha_core/n8452_4 ),
	.I1(\top/processor/sha_core/n8452_5 ),
	.I2(\top/processor/sha_core/n3915_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8452_3 )
);
defparam \top/processor/sha_core/n8452_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8453_s0  (
	.I0(\top/processor/sha_core/n8453_4 ),
	.I1(\top/processor/sha_core/n8453_5 ),
	.I2(\top/processor/sha_core/n3916_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8453_3 )
);
defparam \top/processor/sha_core/n8453_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8454_s0  (
	.I0(\top/processor/sha_core/n8454_4 ),
	.I1(\top/processor/sha_core/n8454_5 ),
	.I2(\top/processor/sha_core/n3917_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8454_3 )
);
defparam \top/processor/sha_core/n8454_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8455_s0  (
	.I0(\top/processor/sha_core/n8455_4 ),
	.I1(\top/processor/sha_core/n8455_5 ),
	.I2(\top/processor/sha_core/n3918_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8455_3 )
);
defparam \top/processor/sha_core/n8455_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8456_s0  (
	.I0(\top/processor/sha_core/n8456_4 ),
	.I1(\top/processor/sha_core/n8456_5 ),
	.I2(\top/processor/sha_core/n3919_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8456_3 )
);
defparam \top/processor/sha_core/n8456_s0 .INIT=16'h77F0;
LUT3 \top/processor/sha_core/n8457_s0  (
	.I0(\top/processor/sha_core/n3920_5 ),
	.I1(\top/processor/sha_core/n8457_4 ),
	.I2(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8457_3 )
);
defparam \top/processor/sha_core/n8457_s0 .INIT=8'h3A;
LUT4 \top/processor/sha_core/n8458_s0  (
	.I0(\top/processor/sha_core/n8458_4 ),
	.I1(\top/processor/sha_core/n8458_5 ),
	.I2(\top/processor/sha_core/n3921_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8458_3 )
);
defparam \top/processor/sha_core/n8458_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8459_s0  (
	.I0(\top/processor/sha_core/n8459_4 ),
	.I1(\top/processor/sha_core/n8459_5 ),
	.I2(\top/processor/sha_core/n3922_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8459_3 )
);
defparam \top/processor/sha_core/n8459_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8460_s0  (
	.I0(\top/processor/sha_core/n8460_4 ),
	.I1(\top/processor/sha_core/n8460_5 ),
	.I2(\top/processor/sha_core/n3923_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8460_3 )
);
defparam \top/processor/sha_core/n8460_s0 .INIT=16'h77F0;
LUT4 \top/processor/sha_core/n8461_s0  (
	.I0(\top/processor/sha_core/n8461_4 ),
	.I1(\top/processor/sha_core/n8461_5 ),
	.I2(\top/processor/sha_core/n3924_5 ),
	.I3(\top/processor/sha_core/n8430_6 ),
	.F(\top/processor/sha_core/n8461_3 )
);
defparam \top/processor/sha_core/n8461_s0 .INIT=16'h77F0;
LUT3 \top/processor/sha_core/n11869_s6  (
	.I0(\top/processor/core_start ),
	.I1(\top/processor/sha_core/state [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11869_11 )
);
defparam \top/processor/sha_core/n11869_s6 .INIT=8'hC2;
LUT3 \top/processor/sha_core/n11872_s5  (
	.I0(\top/processor/sha_core/h7 [31]),
	.I1(\top/processor/sha_core/g [31]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11872_9 )
);
defparam \top/processor/sha_core/n11872_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11873_s5  (
	.I0(\top/processor/sha_core/h7 [30]),
	.I1(\top/processor/sha_core/g [30]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11873_9 )
);
defparam \top/processor/sha_core/n11873_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11874_s5  (
	.I0(\top/processor/sha_core/h7 [29]),
	.I1(\top/processor/sha_core/g [29]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11874_9 )
);
defparam \top/processor/sha_core/n11874_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11875_s5  (
	.I0(\top/processor/sha_core/h7 [28]),
	.I1(\top/processor/sha_core/g [28]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11875_9 )
);
defparam \top/processor/sha_core/n11875_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11876_s5  (
	.I0(\top/processor/sha_core/h7 [27]),
	.I1(\top/processor/sha_core/g [27]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11876_9 )
);
defparam \top/processor/sha_core/n11876_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11877_s5  (
	.I0(\top/processor/sha_core/h7 [26]),
	.I1(\top/processor/sha_core/g [26]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11877_9 )
);
defparam \top/processor/sha_core/n11877_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11878_s5  (
	.I0(\top/processor/sha_core/h7 [25]),
	.I1(\top/processor/sha_core/g [25]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11878_9 )
);
defparam \top/processor/sha_core/n11878_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11879_s5  (
	.I0(\top/processor/sha_core/h7 [24]),
	.I1(\top/processor/sha_core/g [24]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11879_9 )
);
defparam \top/processor/sha_core/n11879_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11880_s5  (
	.I0(\top/processor/sha_core/h7 [23]),
	.I1(\top/processor/sha_core/g [23]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11880_9 )
);
defparam \top/processor/sha_core/n11880_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11881_s5  (
	.I0(\top/processor/sha_core/h7 [22]),
	.I1(\top/processor/sha_core/g [22]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11881_9 )
);
defparam \top/processor/sha_core/n11881_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11882_s5  (
	.I0(\top/processor/sha_core/h7 [21]),
	.I1(\top/processor/sha_core/g [21]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11882_9 )
);
defparam \top/processor/sha_core/n11882_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11883_s5  (
	.I0(\top/processor/sha_core/h7 [20]),
	.I1(\top/processor/sha_core/g [20]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11883_9 )
);
defparam \top/processor/sha_core/n11883_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11884_s5  (
	.I0(\top/processor/sha_core/h7 [19]),
	.I1(\top/processor/sha_core/g [19]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11884_9 )
);
defparam \top/processor/sha_core/n11884_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11885_s5  (
	.I0(\top/processor/sha_core/h7 [18]),
	.I1(\top/processor/sha_core/g [18]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11885_9 )
);
defparam \top/processor/sha_core/n11885_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11886_s5  (
	.I0(\top/processor/sha_core/h7 [17]),
	.I1(\top/processor/sha_core/g [17]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11886_9 )
);
defparam \top/processor/sha_core/n11886_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11887_s5  (
	.I0(\top/processor/sha_core/h7 [16]),
	.I1(\top/processor/sha_core/g [16]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11887_9 )
);
defparam \top/processor/sha_core/n11887_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11888_s5  (
	.I0(\top/processor/sha_core/h7 [15]),
	.I1(\top/processor/sha_core/g [15]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11888_9 )
);
defparam \top/processor/sha_core/n11888_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11889_s5  (
	.I0(\top/processor/sha_core/h7 [14]),
	.I1(\top/processor/sha_core/g [14]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11889_9 )
);
defparam \top/processor/sha_core/n11889_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11890_s5  (
	.I0(\top/processor/sha_core/h7 [13]),
	.I1(\top/processor/sha_core/g [13]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11890_9 )
);
defparam \top/processor/sha_core/n11890_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11891_s5  (
	.I0(\top/processor/sha_core/h7 [12]),
	.I1(\top/processor/sha_core/g [12]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11891_9 )
);
defparam \top/processor/sha_core/n11891_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11892_s5  (
	.I0(\top/processor/sha_core/h7 [11]),
	.I1(\top/processor/sha_core/g [11]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11892_9 )
);
defparam \top/processor/sha_core/n11892_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11893_s5  (
	.I0(\top/processor/sha_core/h7 [10]),
	.I1(\top/processor/sha_core/g [10]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11893_9 )
);
defparam \top/processor/sha_core/n11893_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11894_s5  (
	.I0(\top/processor/sha_core/h7 [9]),
	.I1(\top/processor/sha_core/g [9]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11894_9 )
);
defparam \top/processor/sha_core/n11894_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11895_s5  (
	.I0(\top/processor/sha_core/h7 [8]),
	.I1(\top/processor/sha_core/g [8]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11895_9 )
);
defparam \top/processor/sha_core/n11895_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11896_s5  (
	.I0(\top/processor/sha_core/h7 [7]),
	.I1(\top/processor/sha_core/g [7]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11896_9 )
);
defparam \top/processor/sha_core/n11896_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11897_s5  (
	.I0(\top/processor/sha_core/h7 [6]),
	.I1(\top/processor/sha_core/g [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11897_9 )
);
defparam \top/processor/sha_core/n11897_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11898_s5  (
	.I0(\top/processor/sha_core/h7 [5]),
	.I1(\top/processor/sha_core/g [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11898_9 )
);
defparam \top/processor/sha_core/n11898_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11899_s5  (
	.I0(\top/processor/sha_core/h7 [4]),
	.I1(\top/processor/sha_core/g [4]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11899_9 )
);
defparam \top/processor/sha_core/n11899_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11900_s5  (
	.I0(\top/processor/sha_core/h7 [3]),
	.I1(\top/processor/sha_core/g [3]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11900_9 )
);
defparam \top/processor/sha_core/n11900_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11901_s5  (
	.I0(\top/processor/sha_core/h7 [2]),
	.I1(\top/processor/sha_core/g [2]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11901_9 )
);
defparam \top/processor/sha_core/n11901_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11902_s5  (
	.I0(\top/processor/sha_core/h7 [1]),
	.I1(\top/processor/sha_core/g [1]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11902_9 )
);
defparam \top/processor/sha_core/n11902_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11903_s5  (
	.I0(\top/processor/sha_core/h7 [0]),
	.I1(\top/processor/sha_core/g [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11903_9 )
);
defparam \top/processor/sha_core/n11903_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11904_s5  (
	.I0(\top/processor/sha_core/h6 [31]),
	.I1(\top/processor/sha_core/f [31]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11904_9 )
);
defparam \top/processor/sha_core/n11904_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11905_s5  (
	.I0(\top/processor/sha_core/h6 [30]),
	.I1(\top/processor/sha_core/f [30]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11905_9 )
);
defparam \top/processor/sha_core/n11905_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11906_s5  (
	.I0(\top/processor/sha_core/h6 [29]),
	.I1(\top/processor/sha_core/f [29]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11906_9 )
);
defparam \top/processor/sha_core/n11906_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11907_s5  (
	.I0(\top/processor/sha_core/h6 [28]),
	.I1(\top/processor/sha_core/f [28]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11907_9 )
);
defparam \top/processor/sha_core/n11907_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11908_s5  (
	.I0(\top/processor/sha_core/h6 [27]),
	.I1(\top/processor/sha_core/f [27]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11908_9 )
);
defparam \top/processor/sha_core/n11908_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11909_s5  (
	.I0(\top/processor/sha_core/h6 [26]),
	.I1(\top/processor/sha_core/f [26]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11909_9 )
);
defparam \top/processor/sha_core/n11909_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11910_s5  (
	.I0(\top/processor/sha_core/h6 [25]),
	.I1(\top/processor/sha_core/f [25]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11910_9 )
);
defparam \top/processor/sha_core/n11910_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11911_s5  (
	.I0(\top/processor/sha_core/h6 [24]),
	.I1(\top/processor/sha_core/f [24]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11911_9 )
);
defparam \top/processor/sha_core/n11911_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11912_s5  (
	.I0(\top/processor/sha_core/h6 [23]),
	.I1(\top/processor/sha_core/f [23]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11912_9 )
);
defparam \top/processor/sha_core/n11912_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11913_s5  (
	.I0(\top/processor/sha_core/h6 [22]),
	.I1(\top/processor/sha_core/f [22]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11913_9 )
);
defparam \top/processor/sha_core/n11913_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11914_s5  (
	.I0(\top/processor/sha_core/h6 [21]),
	.I1(\top/processor/sha_core/f [21]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11914_9 )
);
defparam \top/processor/sha_core/n11914_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11915_s5  (
	.I0(\top/processor/sha_core/h6 [20]),
	.I1(\top/processor/sha_core/f [20]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11915_9 )
);
defparam \top/processor/sha_core/n11915_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11916_s5  (
	.I0(\top/processor/sha_core/h6 [19]),
	.I1(\top/processor/sha_core/f [19]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11916_9 )
);
defparam \top/processor/sha_core/n11916_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11917_s5  (
	.I0(\top/processor/sha_core/h6 [18]),
	.I1(\top/processor/sha_core/f [18]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11917_9 )
);
defparam \top/processor/sha_core/n11917_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11918_s5  (
	.I0(\top/processor/sha_core/h6 [17]),
	.I1(\top/processor/sha_core/f [17]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11918_9 )
);
defparam \top/processor/sha_core/n11918_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11919_s5  (
	.I0(\top/processor/sha_core/h6 [16]),
	.I1(\top/processor/sha_core/f [16]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11919_9 )
);
defparam \top/processor/sha_core/n11919_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11920_s5  (
	.I0(\top/processor/sha_core/h6 [15]),
	.I1(\top/processor/sha_core/f [15]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11920_9 )
);
defparam \top/processor/sha_core/n11920_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11921_s5  (
	.I0(\top/processor/sha_core/h6 [14]),
	.I1(\top/processor/sha_core/f [14]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11921_9 )
);
defparam \top/processor/sha_core/n11921_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11922_s5  (
	.I0(\top/processor/sha_core/h6 [13]),
	.I1(\top/processor/sha_core/f [13]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11922_9 )
);
defparam \top/processor/sha_core/n11922_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11923_s5  (
	.I0(\top/processor/sha_core/h6 [12]),
	.I1(\top/processor/sha_core/f [12]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11923_9 )
);
defparam \top/processor/sha_core/n11923_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11924_s5  (
	.I0(\top/processor/sha_core/h6 [11]),
	.I1(\top/processor/sha_core/f [11]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11924_9 )
);
defparam \top/processor/sha_core/n11924_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11925_s5  (
	.I0(\top/processor/sha_core/h6 [10]),
	.I1(\top/processor/sha_core/f [10]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11925_9 )
);
defparam \top/processor/sha_core/n11925_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11926_s5  (
	.I0(\top/processor/sha_core/h6 [9]),
	.I1(\top/processor/sha_core/f [9]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11926_9 )
);
defparam \top/processor/sha_core/n11926_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11927_s5  (
	.I0(\top/processor/sha_core/h6 [8]),
	.I1(\top/processor/sha_core/f [8]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11927_9 )
);
defparam \top/processor/sha_core/n11927_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11928_s5  (
	.I0(\top/processor/sha_core/h6 [7]),
	.I1(\top/processor/sha_core/f [7]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11928_9 )
);
defparam \top/processor/sha_core/n11928_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11929_s5  (
	.I0(\top/processor/sha_core/h6 [6]),
	.I1(\top/processor/sha_core/f [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11929_9 )
);
defparam \top/processor/sha_core/n11929_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11930_s5  (
	.I0(\top/processor/sha_core/h6 [5]),
	.I1(\top/processor/sha_core/f [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11930_9 )
);
defparam \top/processor/sha_core/n11930_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11931_s5  (
	.I0(\top/processor/sha_core/h6 [4]),
	.I1(\top/processor/sha_core/f [4]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11931_9 )
);
defparam \top/processor/sha_core/n11931_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11932_s5  (
	.I0(\top/processor/sha_core/h6 [3]),
	.I1(\top/processor/sha_core/f [3]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11932_9 )
);
defparam \top/processor/sha_core/n11932_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11933_s5  (
	.I0(\top/processor/sha_core/h6 [2]),
	.I1(\top/processor/sha_core/f [2]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11933_9 )
);
defparam \top/processor/sha_core/n11933_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11934_s5  (
	.I0(\top/processor/sha_core/h6 [1]),
	.I1(\top/processor/sha_core/f [1]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11934_9 )
);
defparam \top/processor/sha_core/n11934_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11935_s5  (
	.I0(\top/processor/sha_core/h6 [0]),
	.I1(\top/processor/sha_core/f [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11935_9 )
);
defparam \top/processor/sha_core/n11935_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11936_s5  (
	.I0(\top/processor/sha_core/h5 [31]),
	.I1(\top/processor/sha_core/e [31]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11936_9 )
);
defparam \top/processor/sha_core/n11936_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11937_s5  (
	.I0(\top/processor/sha_core/h5 [30]),
	.I1(\top/processor/sha_core/e [30]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11937_9 )
);
defparam \top/processor/sha_core/n11937_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11938_s5  (
	.I0(\top/processor/sha_core/h5 [29]),
	.I1(\top/processor/sha_core/e [29]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11938_9 )
);
defparam \top/processor/sha_core/n11938_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11939_s5  (
	.I0(\top/processor/sha_core/h5 [28]),
	.I1(\top/processor/sha_core/e [28]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11939_9 )
);
defparam \top/processor/sha_core/n11939_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11940_s5  (
	.I0(\top/processor/sha_core/h5 [27]),
	.I1(\top/processor/sha_core/e [27]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11940_9 )
);
defparam \top/processor/sha_core/n11940_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11941_s5  (
	.I0(\top/processor/sha_core/h5 [26]),
	.I1(\top/processor/sha_core/e [26]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11941_9 )
);
defparam \top/processor/sha_core/n11941_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11942_s5  (
	.I0(\top/processor/sha_core/h5 [25]),
	.I1(\top/processor/sha_core/e [25]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11942_9 )
);
defparam \top/processor/sha_core/n11942_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11943_s5  (
	.I0(\top/processor/sha_core/h5 [24]),
	.I1(\top/processor/sha_core/e [24]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11943_9 )
);
defparam \top/processor/sha_core/n11943_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11944_s5  (
	.I0(\top/processor/sha_core/h5 [23]),
	.I1(\top/processor/sha_core/e [23]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11944_9 )
);
defparam \top/processor/sha_core/n11944_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11945_s5  (
	.I0(\top/processor/sha_core/h5 [22]),
	.I1(\top/processor/sha_core/e [22]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11945_9 )
);
defparam \top/processor/sha_core/n11945_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11946_s5  (
	.I0(\top/processor/sha_core/h5 [21]),
	.I1(\top/processor/sha_core/e [21]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11946_9 )
);
defparam \top/processor/sha_core/n11946_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11947_s5  (
	.I0(\top/processor/sha_core/h5 [20]),
	.I1(\top/processor/sha_core/e [20]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11947_9 )
);
defparam \top/processor/sha_core/n11947_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11948_s5  (
	.I0(\top/processor/sha_core/h5 [19]),
	.I1(\top/processor/sha_core/e [19]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11948_9 )
);
defparam \top/processor/sha_core/n11948_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11949_s5  (
	.I0(\top/processor/sha_core/h5 [18]),
	.I1(\top/processor/sha_core/e [18]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11949_9 )
);
defparam \top/processor/sha_core/n11949_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11950_s5  (
	.I0(\top/processor/sha_core/h5 [17]),
	.I1(\top/processor/sha_core/e [17]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11950_9 )
);
defparam \top/processor/sha_core/n11950_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11951_s5  (
	.I0(\top/processor/sha_core/h5 [16]),
	.I1(\top/processor/sha_core/e [16]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11951_9 )
);
defparam \top/processor/sha_core/n11951_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11952_s5  (
	.I0(\top/processor/sha_core/h5 [15]),
	.I1(\top/processor/sha_core/e [15]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11952_9 )
);
defparam \top/processor/sha_core/n11952_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11953_s5  (
	.I0(\top/processor/sha_core/h5 [14]),
	.I1(\top/processor/sha_core/e [14]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11953_9 )
);
defparam \top/processor/sha_core/n11953_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11954_s5  (
	.I0(\top/processor/sha_core/h5 [13]),
	.I1(\top/processor/sha_core/e [13]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11954_9 )
);
defparam \top/processor/sha_core/n11954_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11955_s5  (
	.I0(\top/processor/sha_core/h5 [12]),
	.I1(\top/processor/sha_core/e [12]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11955_9 )
);
defparam \top/processor/sha_core/n11955_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11956_s5  (
	.I0(\top/processor/sha_core/h5 [11]),
	.I1(\top/processor/sha_core/e [11]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11956_9 )
);
defparam \top/processor/sha_core/n11956_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11957_s5  (
	.I0(\top/processor/sha_core/h5 [10]),
	.I1(\top/processor/sha_core/e [10]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11957_9 )
);
defparam \top/processor/sha_core/n11957_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11958_s5  (
	.I0(\top/processor/sha_core/h5 [9]),
	.I1(\top/processor/sha_core/e [9]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11958_9 )
);
defparam \top/processor/sha_core/n11958_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11959_s5  (
	.I0(\top/processor/sha_core/h5 [8]),
	.I1(\top/processor/sha_core/e [8]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11959_9 )
);
defparam \top/processor/sha_core/n11959_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11960_s5  (
	.I0(\top/processor/sha_core/h5 [7]),
	.I1(\top/processor/sha_core/e [7]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11960_9 )
);
defparam \top/processor/sha_core/n11960_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11961_s5  (
	.I0(\top/processor/sha_core/h5 [6]),
	.I1(\top/processor/sha_core/e [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11961_9 )
);
defparam \top/processor/sha_core/n11961_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11962_s5  (
	.I0(\top/processor/sha_core/h5 [5]),
	.I1(\top/processor/sha_core/e [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11962_9 )
);
defparam \top/processor/sha_core/n11962_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11963_s5  (
	.I0(\top/processor/sha_core/h5 [4]),
	.I1(\top/processor/sha_core/e [4]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11963_9 )
);
defparam \top/processor/sha_core/n11963_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11964_s5  (
	.I0(\top/processor/sha_core/h5 [3]),
	.I1(\top/processor/sha_core/e [3]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11964_9 )
);
defparam \top/processor/sha_core/n11964_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11965_s5  (
	.I0(\top/processor/sha_core/h5 [2]),
	.I1(\top/processor/sha_core/e [2]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11965_9 )
);
defparam \top/processor/sha_core/n11965_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11966_s5  (
	.I0(\top/processor/sha_core/h5 [1]),
	.I1(\top/processor/sha_core/e [1]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11966_9 )
);
defparam \top/processor/sha_core/n11966_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11967_s5  (
	.I0(\top/processor/sha_core/h5 [0]),
	.I1(\top/processor/sha_core/e [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11967_9 )
);
defparam \top/processor/sha_core/n11967_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11968_s5  (
	.I0(\top/processor/sha_core/h4 [31]),
	.I1(\top/processor/sha_core/n10752_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11968_9 )
);
defparam \top/processor/sha_core/n11968_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11969_s5  (
	.I0(\top/processor/sha_core/h4 [30]),
	.I1(\top/processor/sha_core/n10753_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11969_9 )
);
defparam \top/processor/sha_core/n11969_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11970_s5  (
	.I0(\top/processor/sha_core/h4 [29]),
	.I1(\top/processor/sha_core/n10754_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11970_9 )
);
defparam \top/processor/sha_core/n11970_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11971_s5  (
	.I0(\top/processor/sha_core/h4 [28]),
	.I1(\top/processor/sha_core/n10755_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11971_9 )
);
defparam \top/processor/sha_core/n11971_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11972_s5  (
	.I0(\top/processor/sha_core/h4 [27]),
	.I1(\top/processor/sha_core/n10756_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11972_9 )
);
defparam \top/processor/sha_core/n11972_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11973_s5  (
	.I0(\top/processor/sha_core/h4 [26]),
	.I1(\top/processor/sha_core/n10757_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11973_9 )
);
defparam \top/processor/sha_core/n11973_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11974_s5  (
	.I0(\top/processor/sha_core/h4 [25]),
	.I1(\top/processor/sha_core/n10758_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11974_9 )
);
defparam \top/processor/sha_core/n11974_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11975_s5  (
	.I0(\top/processor/sha_core/h4 [24]),
	.I1(\top/processor/sha_core/n10759_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11975_9 )
);
defparam \top/processor/sha_core/n11975_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11976_s5  (
	.I0(\top/processor/sha_core/h4 [23]),
	.I1(\top/processor/sha_core/n10760_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11976_9 )
);
defparam \top/processor/sha_core/n11976_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11977_s5  (
	.I0(\top/processor/sha_core/h4 [22]),
	.I1(\top/processor/sha_core/n10761_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11977_9 )
);
defparam \top/processor/sha_core/n11977_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11978_s5  (
	.I0(\top/processor/sha_core/h4 [21]),
	.I1(\top/processor/sha_core/n10762_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11978_9 )
);
defparam \top/processor/sha_core/n11978_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11979_s5  (
	.I0(\top/processor/sha_core/h4 [20]),
	.I1(\top/processor/sha_core/n10763_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11979_9 )
);
defparam \top/processor/sha_core/n11979_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11980_s5  (
	.I0(\top/processor/sha_core/h4 [19]),
	.I1(\top/processor/sha_core/n10764_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11980_9 )
);
defparam \top/processor/sha_core/n11980_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11981_s5  (
	.I0(\top/processor/sha_core/h4 [18]),
	.I1(\top/processor/sha_core/n10765_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11981_9 )
);
defparam \top/processor/sha_core/n11981_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11982_s5  (
	.I0(\top/processor/sha_core/h4 [17]),
	.I1(\top/processor/sha_core/n10766_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11982_9 )
);
defparam \top/processor/sha_core/n11982_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11983_s5  (
	.I0(\top/processor/sha_core/h4 [16]),
	.I1(\top/processor/sha_core/n10767_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11983_9 )
);
defparam \top/processor/sha_core/n11983_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11984_s5  (
	.I0(\top/processor/sha_core/h4 [15]),
	.I1(\top/processor/sha_core/n10768_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11984_9 )
);
defparam \top/processor/sha_core/n11984_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11985_s5  (
	.I0(\top/processor/sha_core/h4 [14]),
	.I1(\top/processor/sha_core/n10769_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11985_9 )
);
defparam \top/processor/sha_core/n11985_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11986_s5  (
	.I0(\top/processor/sha_core/h4 [13]),
	.I1(\top/processor/sha_core/n10770_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11986_9 )
);
defparam \top/processor/sha_core/n11986_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11987_s5  (
	.I0(\top/processor/sha_core/h4 [12]),
	.I1(\top/processor/sha_core/n10771_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11987_9 )
);
defparam \top/processor/sha_core/n11987_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11988_s5  (
	.I0(\top/processor/sha_core/h4 [11]),
	.I1(\top/processor/sha_core/n10772_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11988_9 )
);
defparam \top/processor/sha_core/n11988_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11989_s5  (
	.I0(\top/processor/sha_core/h4 [10]),
	.I1(\top/processor/sha_core/n10773_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11989_9 )
);
defparam \top/processor/sha_core/n11989_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11990_s5  (
	.I0(\top/processor/sha_core/h4 [9]),
	.I1(\top/processor/sha_core/n10774_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11990_9 )
);
defparam \top/processor/sha_core/n11990_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11991_s5  (
	.I0(\top/processor/sha_core/h4 [8]),
	.I1(\top/processor/sha_core/n10775_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11991_9 )
);
defparam \top/processor/sha_core/n11991_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11992_s5  (
	.I0(\top/processor/sha_core/h4 [7]),
	.I1(\top/processor/sha_core/n10776_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11992_9 )
);
defparam \top/processor/sha_core/n11992_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11993_s5  (
	.I0(\top/processor/sha_core/h4 [6]),
	.I1(\top/processor/sha_core/n10777_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11993_9 )
);
defparam \top/processor/sha_core/n11993_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11994_s5  (
	.I0(\top/processor/sha_core/h4 [5]),
	.I1(\top/processor/sha_core/n10778_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11994_9 )
);
defparam \top/processor/sha_core/n11994_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11995_s5  (
	.I0(\top/processor/sha_core/h4 [4]),
	.I1(\top/processor/sha_core/n10779_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11995_9 )
);
defparam \top/processor/sha_core/n11995_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11996_s5  (
	.I0(\top/processor/sha_core/h4 [3]),
	.I1(\top/processor/sha_core/n10780_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11996_9 )
);
defparam \top/processor/sha_core/n11996_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11997_s5  (
	.I0(\top/processor/sha_core/h4 [2]),
	.I1(\top/processor/sha_core/n10781_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11997_9 )
);
defparam \top/processor/sha_core/n11997_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11998_s5  (
	.I0(\top/processor/sha_core/h4 [1]),
	.I1(\top/processor/sha_core/n10782_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11998_9 )
);
defparam \top/processor/sha_core/n11998_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n11999_s5  (
	.I0(\top/processor/sha_core/h4 [0]),
	.I1(\top/processor/sha_core/n10783_11 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11999_9 )
);
defparam \top/processor/sha_core/n11999_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12000_s5  (
	.I0(\top/processor/sha_core/h3 [31]),
	.I1(\top/processor/sha_core/c [31]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12000_9 )
);
defparam \top/processor/sha_core/n12000_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12001_s5  (
	.I0(\top/processor/sha_core/h3 [30]),
	.I1(\top/processor/sha_core/c [30]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12001_9 )
);
defparam \top/processor/sha_core/n12001_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12002_s5  (
	.I0(\top/processor/sha_core/h3 [29]),
	.I1(\top/processor/sha_core/c [29]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12002_9 )
);
defparam \top/processor/sha_core/n12002_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12003_s5  (
	.I0(\top/processor/sha_core/h3 [28]),
	.I1(\top/processor/sha_core/c [28]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12003_9 )
);
defparam \top/processor/sha_core/n12003_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12004_s5  (
	.I0(\top/processor/sha_core/h3 [27]),
	.I1(\top/processor/sha_core/c [27]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12004_9 )
);
defparam \top/processor/sha_core/n12004_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12005_s5  (
	.I0(\top/processor/sha_core/h3 [26]),
	.I1(\top/processor/sha_core/c [26]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12005_9 )
);
defparam \top/processor/sha_core/n12005_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12006_s5  (
	.I0(\top/processor/sha_core/h3 [25]),
	.I1(\top/processor/sha_core/c [25]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12006_9 )
);
defparam \top/processor/sha_core/n12006_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12007_s5  (
	.I0(\top/processor/sha_core/h3 [24]),
	.I1(\top/processor/sha_core/c [24]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12007_9 )
);
defparam \top/processor/sha_core/n12007_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12008_s5  (
	.I0(\top/processor/sha_core/h3 [23]),
	.I1(\top/processor/sha_core/c [23]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12008_9 )
);
defparam \top/processor/sha_core/n12008_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12009_s5  (
	.I0(\top/processor/sha_core/h3 [22]),
	.I1(\top/processor/sha_core/c [22]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12009_9 )
);
defparam \top/processor/sha_core/n12009_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12010_s5  (
	.I0(\top/processor/sha_core/h3 [21]),
	.I1(\top/processor/sha_core/c [21]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12010_9 )
);
defparam \top/processor/sha_core/n12010_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12011_s5  (
	.I0(\top/processor/sha_core/h3 [20]),
	.I1(\top/processor/sha_core/c [20]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12011_9 )
);
defparam \top/processor/sha_core/n12011_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12012_s5  (
	.I0(\top/processor/sha_core/h3 [19]),
	.I1(\top/processor/sha_core/c [19]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12012_9 )
);
defparam \top/processor/sha_core/n12012_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12013_s5  (
	.I0(\top/processor/sha_core/h3 [18]),
	.I1(\top/processor/sha_core/c [18]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12013_9 )
);
defparam \top/processor/sha_core/n12013_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12014_s5  (
	.I0(\top/processor/sha_core/h3 [17]),
	.I1(\top/processor/sha_core/c [17]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12014_9 )
);
defparam \top/processor/sha_core/n12014_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12015_s5  (
	.I0(\top/processor/sha_core/h3 [16]),
	.I1(\top/processor/sha_core/c [16]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12015_9 )
);
defparam \top/processor/sha_core/n12015_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12016_s5  (
	.I0(\top/processor/sha_core/h3 [15]),
	.I1(\top/processor/sha_core/c [15]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12016_9 )
);
defparam \top/processor/sha_core/n12016_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12017_s5  (
	.I0(\top/processor/sha_core/h3 [14]),
	.I1(\top/processor/sha_core/c [14]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12017_9 )
);
defparam \top/processor/sha_core/n12017_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12018_s5  (
	.I0(\top/processor/sha_core/h3 [13]),
	.I1(\top/processor/sha_core/c [13]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12018_9 )
);
defparam \top/processor/sha_core/n12018_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12019_s5  (
	.I0(\top/processor/sha_core/h3 [12]),
	.I1(\top/processor/sha_core/c [12]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12019_9 )
);
defparam \top/processor/sha_core/n12019_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12020_s5  (
	.I0(\top/processor/sha_core/h3 [11]),
	.I1(\top/processor/sha_core/c [11]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12020_9 )
);
defparam \top/processor/sha_core/n12020_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12021_s5  (
	.I0(\top/processor/sha_core/h3 [10]),
	.I1(\top/processor/sha_core/c [10]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12021_9 )
);
defparam \top/processor/sha_core/n12021_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12022_s5  (
	.I0(\top/processor/sha_core/h3 [9]),
	.I1(\top/processor/sha_core/c [9]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12022_9 )
);
defparam \top/processor/sha_core/n12022_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12023_s5  (
	.I0(\top/processor/sha_core/h3 [8]),
	.I1(\top/processor/sha_core/c [8]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12023_9 )
);
defparam \top/processor/sha_core/n12023_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12024_s5  (
	.I0(\top/processor/sha_core/h3 [7]),
	.I1(\top/processor/sha_core/c [7]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12024_9 )
);
defparam \top/processor/sha_core/n12024_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12025_s5  (
	.I0(\top/processor/sha_core/h3 [6]),
	.I1(\top/processor/sha_core/c [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12025_9 )
);
defparam \top/processor/sha_core/n12025_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12026_s5  (
	.I0(\top/processor/sha_core/h3 [5]),
	.I1(\top/processor/sha_core/c [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12026_9 )
);
defparam \top/processor/sha_core/n12026_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12027_s5  (
	.I0(\top/processor/sha_core/h3 [4]),
	.I1(\top/processor/sha_core/c [4]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12027_9 )
);
defparam \top/processor/sha_core/n12027_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12028_s5  (
	.I0(\top/processor/sha_core/h3 [3]),
	.I1(\top/processor/sha_core/c [3]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12028_9 )
);
defparam \top/processor/sha_core/n12028_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12029_s5  (
	.I0(\top/processor/sha_core/h3 [2]),
	.I1(\top/processor/sha_core/c [2]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12029_9 )
);
defparam \top/processor/sha_core/n12029_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12030_s5  (
	.I0(\top/processor/sha_core/h3 [1]),
	.I1(\top/processor/sha_core/c [1]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12030_9 )
);
defparam \top/processor/sha_core/n12030_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12031_s5  (
	.I0(\top/processor/sha_core/h3 [0]),
	.I1(\top/processor/sha_core/c [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12031_9 )
);
defparam \top/processor/sha_core/n12031_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12032_s5  (
	.I0(\top/processor/sha_core/h2 [31]),
	.I1(\top/processor/sha_core/b [31]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12032_9 )
);
defparam \top/processor/sha_core/n12032_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12033_s5  (
	.I0(\top/processor/sha_core/h2 [30]),
	.I1(\top/processor/sha_core/b [30]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12033_9 )
);
defparam \top/processor/sha_core/n12033_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12034_s5  (
	.I0(\top/processor/sha_core/h2 [29]),
	.I1(\top/processor/sha_core/b [29]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12034_9 )
);
defparam \top/processor/sha_core/n12034_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12035_s5  (
	.I0(\top/processor/sha_core/h2 [28]),
	.I1(\top/processor/sha_core/b [28]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12035_9 )
);
defparam \top/processor/sha_core/n12035_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12036_s5  (
	.I0(\top/processor/sha_core/h2 [27]),
	.I1(\top/processor/sha_core/b [27]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12036_9 )
);
defparam \top/processor/sha_core/n12036_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12037_s5  (
	.I0(\top/processor/sha_core/h2 [26]),
	.I1(\top/processor/sha_core/b [26]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12037_9 )
);
defparam \top/processor/sha_core/n12037_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12038_s5  (
	.I0(\top/processor/sha_core/h2 [25]),
	.I1(\top/processor/sha_core/b [25]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12038_9 )
);
defparam \top/processor/sha_core/n12038_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12039_s5  (
	.I0(\top/processor/sha_core/h2 [24]),
	.I1(\top/processor/sha_core/b [24]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12039_9 )
);
defparam \top/processor/sha_core/n12039_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12040_s5  (
	.I0(\top/processor/sha_core/h2 [23]),
	.I1(\top/processor/sha_core/b [23]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12040_9 )
);
defparam \top/processor/sha_core/n12040_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12041_s5  (
	.I0(\top/processor/sha_core/h2 [22]),
	.I1(\top/processor/sha_core/b [22]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12041_9 )
);
defparam \top/processor/sha_core/n12041_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12042_s5  (
	.I0(\top/processor/sha_core/h2 [21]),
	.I1(\top/processor/sha_core/b [21]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12042_9 )
);
defparam \top/processor/sha_core/n12042_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12043_s5  (
	.I0(\top/processor/sha_core/h2 [20]),
	.I1(\top/processor/sha_core/b [20]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12043_9 )
);
defparam \top/processor/sha_core/n12043_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12044_s5  (
	.I0(\top/processor/sha_core/h2 [19]),
	.I1(\top/processor/sha_core/b [19]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12044_9 )
);
defparam \top/processor/sha_core/n12044_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12045_s5  (
	.I0(\top/processor/sha_core/h2 [18]),
	.I1(\top/processor/sha_core/b [18]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12045_9 )
);
defparam \top/processor/sha_core/n12045_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12046_s5  (
	.I0(\top/processor/sha_core/h2 [17]),
	.I1(\top/processor/sha_core/b [17]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12046_9 )
);
defparam \top/processor/sha_core/n12046_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12047_s5  (
	.I0(\top/processor/sha_core/h2 [16]),
	.I1(\top/processor/sha_core/b [16]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12047_9 )
);
defparam \top/processor/sha_core/n12047_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12048_s5  (
	.I0(\top/processor/sha_core/h2 [15]),
	.I1(\top/processor/sha_core/b [15]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12048_9 )
);
defparam \top/processor/sha_core/n12048_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12049_s5  (
	.I0(\top/processor/sha_core/h2 [14]),
	.I1(\top/processor/sha_core/b [14]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12049_9 )
);
defparam \top/processor/sha_core/n12049_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12050_s5  (
	.I0(\top/processor/sha_core/h2 [13]),
	.I1(\top/processor/sha_core/b [13]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12050_9 )
);
defparam \top/processor/sha_core/n12050_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12051_s5  (
	.I0(\top/processor/sha_core/h2 [12]),
	.I1(\top/processor/sha_core/b [12]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12051_9 )
);
defparam \top/processor/sha_core/n12051_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12052_s5  (
	.I0(\top/processor/sha_core/h2 [11]),
	.I1(\top/processor/sha_core/b [11]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12052_9 )
);
defparam \top/processor/sha_core/n12052_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12053_s5  (
	.I0(\top/processor/sha_core/h2 [10]),
	.I1(\top/processor/sha_core/b [10]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12053_9 )
);
defparam \top/processor/sha_core/n12053_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12054_s5  (
	.I0(\top/processor/sha_core/h2 [9]),
	.I1(\top/processor/sha_core/b [9]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12054_9 )
);
defparam \top/processor/sha_core/n12054_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12055_s5  (
	.I0(\top/processor/sha_core/h2 [8]),
	.I1(\top/processor/sha_core/b [8]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12055_9 )
);
defparam \top/processor/sha_core/n12055_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12056_s5  (
	.I0(\top/processor/sha_core/h2 [7]),
	.I1(\top/processor/sha_core/b [7]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12056_9 )
);
defparam \top/processor/sha_core/n12056_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12057_s5  (
	.I0(\top/processor/sha_core/h2 [6]),
	.I1(\top/processor/sha_core/b [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12057_9 )
);
defparam \top/processor/sha_core/n12057_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12058_s5  (
	.I0(\top/processor/sha_core/h2 [5]),
	.I1(\top/processor/sha_core/b [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12058_9 )
);
defparam \top/processor/sha_core/n12058_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12059_s5  (
	.I0(\top/processor/sha_core/h2 [4]),
	.I1(\top/processor/sha_core/b [4]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12059_9 )
);
defparam \top/processor/sha_core/n12059_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12060_s5  (
	.I0(\top/processor/sha_core/h2 [3]),
	.I1(\top/processor/sha_core/b [3]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12060_9 )
);
defparam \top/processor/sha_core/n12060_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12061_s5  (
	.I0(\top/processor/sha_core/h2 [2]),
	.I1(\top/processor/sha_core/b [2]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12061_9 )
);
defparam \top/processor/sha_core/n12061_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12062_s5  (
	.I0(\top/processor/sha_core/h2 [1]),
	.I1(\top/processor/sha_core/b [1]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12062_9 )
);
defparam \top/processor/sha_core/n12062_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12063_s5  (
	.I0(\top/processor/sha_core/h2 [0]),
	.I1(\top/processor/sha_core/b [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12063_9 )
);
defparam \top/processor/sha_core/n12063_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12064_s5  (
	.I0(\top/processor/sha_core/h1 [31]),
	.I1(\top/processor/sha_core/a [31]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12064_9 )
);
defparam \top/processor/sha_core/n12064_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12065_s5  (
	.I0(\top/processor/sha_core/h1 [30]),
	.I1(\top/processor/sha_core/a [30]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12065_9 )
);
defparam \top/processor/sha_core/n12065_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12066_s5  (
	.I0(\top/processor/sha_core/h1 [29]),
	.I1(\top/processor/sha_core/a [29]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12066_9 )
);
defparam \top/processor/sha_core/n12066_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12067_s5  (
	.I0(\top/processor/sha_core/h1 [28]),
	.I1(\top/processor/sha_core/a [28]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12067_9 )
);
defparam \top/processor/sha_core/n12067_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12068_s5  (
	.I0(\top/processor/sha_core/h1 [27]),
	.I1(\top/processor/sha_core/a [27]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12068_9 )
);
defparam \top/processor/sha_core/n12068_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12069_s5  (
	.I0(\top/processor/sha_core/h1 [26]),
	.I1(\top/processor/sha_core/a [26]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12069_9 )
);
defparam \top/processor/sha_core/n12069_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12070_s5  (
	.I0(\top/processor/sha_core/h1 [25]),
	.I1(\top/processor/sha_core/a [25]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12070_9 )
);
defparam \top/processor/sha_core/n12070_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12071_s5  (
	.I0(\top/processor/sha_core/h1 [24]),
	.I1(\top/processor/sha_core/a [24]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12071_9 )
);
defparam \top/processor/sha_core/n12071_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12072_s5  (
	.I0(\top/processor/sha_core/h1 [23]),
	.I1(\top/processor/sha_core/a [23]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12072_9 )
);
defparam \top/processor/sha_core/n12072_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12073_s5  (
	.I0(\top/processor/sha_core/h1 [22]),
	.I1(\top/processor/sha_core/a [22]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12073_9 )
);
defparam \top/processor/sha_core/n12073_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12074_s5  (
	.I0(\top/processor/sha_core/h1 [21]),
	.I1(\top/processor/sha_core/a [21]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12074_9 )
);
defparam \top/processor/sha_core/n12074_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12075_s5  (
	.I0(\top/processor/sha_core/h1 [20]),
	.I1(\top/processor/sha_core/a [20]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12075_9 )
);
defparam \top/processor/sha_core/n12075_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12076_s5  (
	.I0(\top/processor/sha_core/h1 [19]),
	.I1(\top/processor/sha_core/a [19]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12076_9 )
);
defparam \top/processor/sha_core/n12076_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12077_s5  (
	.I0(\top/processor/sha_core/h1 [18]),
	.I1(\top/processor/sha_core/a [18]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12077_9 )
);
defparam \top/processor/sha_core/n12077_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12078_s5  (
	.I0(\top/processor/sha_core/h1 [17]),
	.I1(\top/processor/sha_core/a [17]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12078_9 )
);
defparam \top/processor/sha_core/n12078_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12079_s5  (
	.I0(\top/processor/sha_core/h1 [16]),
	.I1(\top/processor/sha_core/a [16]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12079_9 )
);
defparam \top/processor/sha_core/n12079_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12080_s5  (
	.I0(\top/processor/sha_core/h1 [15]),
	.I1(\top/processor/sha_core/a [15]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12080_9 )
);
defparam \top/processor/sha_core/n12080_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12081_s5  (
	.I0(\top/processor/sha_core/h1 [14]),
	.I1(\top/processor/sha_core/a [14]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12081_9 )
);
defparam \top/processor/sha_core/n12081_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12082_s5  (
	.I0(\top/processor/sha_core/h1 [13]),
	.I1(\top/processor/sha_core/a [13]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12082_9 )
);
defparam \top/processor/sha_core/n12082_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12083_s5  (
	.I0(\top/processor/sha_core/h1 [12]),
	.I1(\top/processor/sha_core/a [12]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12083_9 )
);
defparam \top/processor/sha_core/n12083_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12084_s5  (
	.I0(\top/processor/sha_core/h1 [11]),
	.I1(\top/processor/sha_core/a [11]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12084_9 )
);
defparam \top/processor/sha_core/n12084_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12085_s5  (
	.I0(\top/processor/sha_core/h1 [10]),
	.I1(\top/processor/sha_core/a [10]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12085_9 )
);
defparam \top/processor/sha_core/n12085_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12086_s5  (
	.I0(\top/processor/sha_core/h1 [9]),
	.I1(\top/processor/sha_core/a [9]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12086_9 )
);
defparam \top/processor/sha_core/n12086_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12087_s5  (
	.I0(\top/processor/sha_core/h1 [8]),
	.I1(\top/processor/sha_core/a [8]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12087_9 )
);
defparam \top/processor/sha_core/n12087_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12088_s5  (
	.I0(\top/processor/sha_core/h1 [7]),
	.I1(\top/processor/sha_core/a [7]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12088_9 )
);
defparam \top/processor/sha_core/n12088_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12089_s5  (
	.I0(\top/processor/sha_core/h1 [6]),
	.I1(\top/processor/sha_core/a [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12089_9 )
);
defparam \top/processor/sha_core/n12089_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12090_s5  (
	.I0(\top/processor/sha_core/h1 [5]),
	.I1(\top/processor/sha_core/a [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12090_9 )
);
defparam \top/processor/sha_core/n12090_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12091_s5  (
	.I0(\top/processor/sha_core/h1 [4]),
	.I1(\top/processor/sha_core/a [4]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12091_9 )
);
defparam \top/processor/sha_core/n12091_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12092_s5  (
	.I0(\top/processor/sha_core/h1 [3]),
	.I1(\top/processor/sha_core/a [3]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12092_9 )
);
defparam \top/processor/sha_core/n12092_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12093_s5  (
	.I0(\top/processor/sha_core/h1 [2]),
	.I1(\top/processor/sha_core/a [2]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12093_9 )
);
defparam \top/processor/sha_core/n12093_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12094_s5  (
	.I0(\top/processor/sha_core/h1 [1]),
	.I1(\top/processor/sha_core/a [1]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12094_9 )
);
defparam \top/processor/sha_core/n12094_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12095_s5  (
	.I0(\top/processor/sha_core/h1 [0]),
	.I1(\top/processor/sha_core/a [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12095_9 )
);
defparam \top/processor/sha_core/n12095_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12096_s5  (
	.I0(\top/processor/sha_core/h0 [31]),
	.I1(\top/processor/sha_core/n10785_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12096_9 )
);
defparam \top/processor/sha_core/n12096_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12097_s5  (
	.I0(\top/processor/sha_core/h0 [30]),
	.I1(\top/processor/sha_core/n10786_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12097_9 )
);
defparam \top/processor/sha_core/n12097_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12098_s5  (
	.I0(\top/processor/sha_core/h0 [29]),
	.I1(\top/processor/sha_core/n10787_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12098_9 )
);
defparam \top/processor/sha_core/n12098_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12099_s5  (
	.I0(\top/processor/sha_core/h0 [28]),
	.I1(\top/processor/sha_core/n10788_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12099_9 )
);
defparam \top/processor/sha_core/n12099_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12100_s5  (
	.I0(\top/processor/sha_core/h0 [27]),
	.I1(\top/processor/sha_core/n10789_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12100_9 )
);
defparam \top/processor/sha_core/n12100_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12101_s5  (
	.I0(\top/processor/sha_core/h0 [26]),
	.I1(\top/processor/sha_core/n10790_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12101_9 )
);
defparam \top/processor/sha_core/n12101_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12102_s5  (
	.I0(\top/processor/sha_core/h0 [25]),
	.I1(\top/processor/sha_core/n10791_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12102_9 )
);
defparam \top/processor/sha_core/n12102_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12103_s5  (
	.I0(\top/processor/sha_core/h0 [24]),
	.I1(\top/processor/sha_core/n10792_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12103_9 )
);
defparam \top/processor/sha_core/n12103_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12104_s5  (
	.I0(\top/processor/sha_core/h0 [23]),
	.I1(\top/processor/sha_core/n10793_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12104_9 )
);
defparam \top/processor/sha_core/n12104_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12105_s5  (
	.I0(\top/processor/sha_core/h0 [22]),
	.I1(\top/processor/sha_core/n10794_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12105_9 )
);
defparam \top/processor/sha_core/n12105_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12106_s5  (
	.I0(\top/processor/sha_core/h0 [21]),
	.I1(\top/processor/sha_core/n10795_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12106_9 )
);
defparam \top/processor/sha_core/n12106_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12107_s5  (
	.I0(\top/processor/sha_core/h0 [20]),
	.I1(\top/processor/sha_core/n10796_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12107_9 )
);
defparam \top/processor/sha_core/n12107_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12108_s5  (
	.I0(\top/processor/sha_core/h0 [19]),
	.I1(\top/processor/sha_core/n10797_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12108_9 )
);
defparam \top/processor/sha_core/n12108_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12109_s5  (
	.I0(\top/processor/sha_core/h0 [18]),
	.I1(\top/processor/sha_core/n10798_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12109_9 )
);
defparam \top/processor/sha_core/n12109_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12110_s5  (
	.I0(\top/processor/sha_core/h0 [17]),
	.I1(\top/processor/sha_core/n10799_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12110_9 )
);
defparam \top/processor/sha_core/n12110_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12111_s5  (
	.I0(\top/processor/sha_core/h0 [16]),
	.I1(\top/processor/sha_core/n10800_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12111_9 )
);
defparam \top/processor/sha_core/n12111_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12112_s5  (
	.I0(\top/processor/sha_core/h0 [15]),
	.I1(\top/processor/sha_core/n10801_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12112_9 )
);
defparam \top/processor/sha_core/n12112_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12113_s5  (
	.I0(\top/processor/sha_core/h0 [14]),
	.I1(\top/processor/sha_core/n10802_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12113_9 )
);
defparam \top/processor/sha_core/n12113_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12114_s5  (
	.I0(\top/processor/sha_core/h0 [13]),
	.I1(\top/processor/sha_core/n10803_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12114_9 )
);
defparam \top/processor/sha_core/n12114_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12115_s5  (
	.I0(\top/processor/sha_core/h0 [12]),
	.I1(\top/processor/sha_core/n10804_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12115_9 )
);
defparam \top/processor/sha_core/n12115_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12116_s5  (
	.I0(\top/processor/sha_core/h0 [11]),
	.I1(\top/processor/sha_core/n10805_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12116_9 )
);
defparam \top/processor/sha_core/n12116_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12117_s5  (
	.I0(\top/processor/sha_core/h0 [10]),
	.I1(\top/processor/sha_core/n10806_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12117_9 )
);
defparam \top/processor/sha_core/n12117_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12118_s5  (
	.I0(\top/processor/sha_core/h0 [9]),
	.I1(\top/processor/sha_core/n10807_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12118_9 )
);
defparam \top/processor/sha_core/n12118_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12119_s5  (
	.I0(\top/processor/sha_core/h0 [8]),
	.I1(\top/processor/sha_core/n10808_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12119_9 )
);
defparam \top/processor/sha_core/n12119_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12120_s5  (
	.I0(\top/processor/sha_core/h0 [7]),
	.I1(\top/processor/sha_core/n10809_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12120_9 )
);
defparam \top/processor/sha_core/n12120_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12121_s5  (
	.I0(\top/processor/sha_core/h0 [6]),
	.I1(\top/processor/sha_core/n10810_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12121_9 )
);
defparam \top/processor/sha_core/n12121_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12122_s5  (
	.I0(\top/processor/sha_core/h0 [5]),
	.I1(\top/processor/sha_core/n10811_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12122_9 )
);
defparam \top/processor/sha_core/n12122_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12123_s5  (
	.I0(\top/processor/sha_core/h0 [4]),
	.I1(\top/processor/sha_core/n10812_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12123_9 )
);
defparam \top/processor/sha_core/n12123_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12124_s5  (
	.I0(\top/processor/sha_core/h0 [3]),
	.I1(\top/processor/sha_core/n10813_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12124_9 )
);
defparam \top/processor/sha_core/n12124_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12125_s5  (
	.I0(\top/processor/sha_core/h0 [2]),
	.I1(\top/processor/sha_core/n10814_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12125_9 )
);
defparam \top/processor/sha_core/n12125_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12126_s5  (
	.I0(\top/processor/sha_core/h0 [1]),
	.I1(\top/processor/sha_core/n10815_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12126_9 )
);
defparam \top/processor/sha_core/n12126_s5 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n12127_s5  (
	.I0(\top/processor/sha_core/h0 [0]),
	.I1(\top/processor/sha_core/n10816_13 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12127_9 )
);
defparam \top/processor/sha_core/n12127_s5 .INIT=8'hCA;
LUT4 \top/processor/sha_core/n12135_s6  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [255]),
	.I2(\top/processor/sha_core/n10826_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12135_10 )
);
defparam \top/processor/sha_core/n12135_s6 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12136_s5  (
	.I0(\top/processor/core_hash_init [254]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10827_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12136_9 )
);
defparam \top/processor/sha_core/n12136_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12137_s5  (
	.I0(\top/processor/core_hash_init [253]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10828_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12137_9 )
);
defparam \top/processor/sha_core/n12137_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12138_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [252]),
	.I2(\top/processor/sha_core/n10829_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12138_9 )
);
defparam \top/processor/sha_core/n12138_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12139_s5  (
	.I0(\top/processor/core_hash_init [251]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10830_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12139_9 )
);
defparam \top/processor/sha_core/n12139_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12140_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [250]),
	.I2(\top/processor/sha_core/n10831_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12140_9 )
);
defparam \top/processor/sha_core/n12140_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12141_s5  (
	.I0(\top/processor/core_hash_init [249]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10832_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12141_9 )
);
defparam \top/processor/sha_core/n12141_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12142_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [248]),
	.I2(\top/processor/sha_core/n10833_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12142_9 )
);
defparam \top/processor/sha_core/n12142_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12143_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [247]),
	.I2(\top/processor/sha_core/n10834_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12143_9 )
);
defparam \top/processor/sha_core/n12143_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12144_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [246]),
	.I2(\top/processor/sha_core/n10835_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12144_9 )
);
defparam \top/processor/sha_core/n12144_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12145_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [245]),
	.I2(\top/processor/sha_core/n10836_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12145_9 )
);
defparam \top/processor/sha_core/n12145_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12146_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [244]),
	.I2(\top/processor/sha_core/n10837_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12146_9 )
);
defparam \top/processor/sha_core/n12146_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12147_s5  (
	.I0(\top/processor/core_hash_init [243]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10838_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12147_9 )
);
defparam \top/processor/sha_core/n12147_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12148_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [242]),
	.I2(\top/processor/sha_core/n10839_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12148_9 )
);
defparam \top/processor/sha_core/n12148_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12149_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [241]),
	.I2(\top/processor/sha_core/n10840_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12149_9 )
);
defparam \top/processor/sha_core/n12149_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12150_s5  (
	.I0(\top/processor/core_hash_init [240]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10841_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12150_9 )
);
defparam \top/processor/sha_core/n12150_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12151_s5  (
	.I0(\top/processor/core_hash_init [239]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10842_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12151_9 )
);
defparam \top/processor/sha_core/n12151_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12152_s5  (
	.I0(\top/processor/core_hash_init [238]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10843_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12152_9 )
);
defparam \top/processor/sha_core/n12152_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12153_s5  (
	.I0(\top/processor/core_hash_init [237]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10844_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12153_9 )
);
defparam \top/processor/sha_core/n12153_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12154_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [236]),
	.I2(\top/processor/sha_core/n10845_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12154_9 )
);
defparam \top/processor/sha_core/n12154_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12155_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [235]),
	.I2(\top/processor/sha_core/n10846_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12155_9 )
);
defparam \top/processor/sha_core/n12155_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12156_s5  (
	.I0(\top/processor/core_hash_init [234]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10847_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12156_9 )
);
defparam \top/processor/sha_core/n12156_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12157_s5  (
	.I0(\top/processor/core_hash_init [233]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10848_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12157_9 )
);
defparam \top/processor/sha_core/n12157_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12158_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [232]),
	.I2(\top/processor/sha_core/n10849_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12158_9 )
);
defparam \top/processor/sha_core/n12158_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12159_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [231]),
	.I2(\top/processor/sha_core/n10850_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12159_9 )
);
defparam \top/processor/sha_core/n12159_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12160_s5  (
	.I0(\top/processor/core_hash_init [230]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10851_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12160_9 )
);
defparam \top/processor/sha_core/n12160_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12161_s5  (
	.I0(\top/processor/core_hash_init [229]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10852_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12161_9 )
);
defparam \top/processor/sha_core/n12161_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12162_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [228]),
	.I2(\top/processor/sha_core/n10853_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12162_9 )
);
defparam \top/processor/sha_core/n12162_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12163_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [227]),
	.I2(\top/processor/sha_core/n10854_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12163_9 )
);
defparam \top/processor/sha_core/n12163_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12164_s5  (
	.I0(\top/processor/core_hash_init [226]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10855_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12164_9 )
);
defparam \top/processor/sha_core/n12164_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12165_s5  (
	.I0(\top/processor/core_hash_init [225]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10856_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12165_9 )
);
defparam \top/processor/sha_core/n12165_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12166_s5  (
	.I0(\top/processor/core_hash_init [224]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10857_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12166_9 )
);
defparam \top/processor/sha_core/n12166_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12167_s5  (
	.I0(\top/processor/core_hash_init [223]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10859_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12167_9 )
);
defparam \top/processor/sha_core/n12167_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12168_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [222]),
	.I2(\top/processor/sha_core/n10860_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12168_9 )
);
defparam \top/processor/sha_core/n12168_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12169_s5  (
	.I0(\top/processor/core_hash_init [221]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10861_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12169_9 )
);
defparam \top/processor/sha_core/n12169_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12170_s5  (
	.I0(\top/processor/core_hash_init [220]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10862_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12170_9 )
);
defparam \top/processor/sha_core/n12170_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12171_s5  (
	.I0(\top/processor/core_hash_init [219]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10863_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12171_9 )
);
defparam \top/processor/sha_core/n12171_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12172_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [218]),
	.I2(\top/processor/sha_core/n10864_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12172_9 )
);
defparam \top/processor/sha_core/n12172_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12173_s5  (
	.I0(\top/processor/core_hash_init [217]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10865_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12173_9 )
);
defparam \top/processor/sha_core/n12173_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12174_s5  (
	.I0(\top/processor/core_hash_init [216]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10866_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12174_9 )
);
defparam \top/processor/sha_core/n12174_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12175_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [215]),
	.I2(\top/processor/sha_core/n10867_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12175_9 )
);
defparam \top/processor/sha_core/n12175_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12176_s5  (
	.I0(\top/processor/core_hash_init [214]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10868_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12176_9 )
);
defparam \top/processor/sha_core/n12176_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12177_s5  (
	.I0(\top/processor/core_hash_init [213]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10869_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12177_9 )
);
defparam \top/processor/sha_core/n12177_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12178_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [212]),
	.I2(\top/processor/sha_core/n10870_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12178_9 )
);
defparam \top/processor/sha_core/n12178_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12179_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [211]),
	.I2(\top/processor/sha_core/n10871_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12179_9 )
);
defparam \top/processor/sha_core/n12179_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12180_s5  (
	.I0(\top/processor/core_hash_init [210]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10872_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12180_9 )
);
defparam \top/processor/sha_core/n12180_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12181_s5  (
	.I0(\top/processor/core_hash_init [209]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10873_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12181_9 )
);
defparam \top/processor/sha_core/n12181_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12182_s5  (
	.I0(\top/processor/core_hash_init [208]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10874_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12182_9 )
);
defparam \top/processor/sha_core/n12182_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12183_s5  (
	.I0(\top/processor/core_hash_init [207]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10875_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12183_9 )
);
defparam \top/processor/sha_core/n12183_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12184_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [206]),
	.I2(\top/processor/sha_core/n10876_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12184_9 )
);
defparam \top/processor/sha_core/n12184_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12185_s5  (
	.I0(\top/processor/core_hash_init [205]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10877_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12185_9 )
);
defparam \top/processor/sha_core/n12185_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12186_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [204]),
	.I2(\top/processor/sha_core/n10878_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12186_9 )
);
defparam \top/processor/sha_core/n12186_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12187_s5  (
	.I0(\top/processor/core_hash_init [203]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10879_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12187_9 )
);
defparam \top/processor/sha_core/n12187_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12188_s5  (
	.I0(\top/processor/core_hash_init [202]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10880_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12188_9 )
);
defparam \top/processor/sha_core/n12188_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12189_s5  (
	.I0(\top/processor/core_hash_init [201]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10881_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12189_9 )
);
defparam \top/processor/sha_core/n12189_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12190_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [200]),
	.I2(\top/processor/sha_core/n10882_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12190_9 )
);
defparam \top/processor/sha_core/n12190_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12191_s5  (
	.I0(\top/processor/core_hash_init [199]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10883_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12191_9 )
);
defparam \top/processor/sha_core/n12191_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12192_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [198]),
	.I2(\top/processor/sha_core/n10884_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12192_9 )
);
defparam \top/processor/sha_core/n12192_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12193_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [197]),
	.I2(\top/processor/sha_core/n10885_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12193_9 )
);
defparam \top/processor/sha_core/n12193_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12194_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [196]),
	.I2(\top/processor/sha_core/n10886_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12194_9 )
);
defparam \top/processor/sha_core/n12194_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12195_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [195]),
	.I2(\top/processor/sha_core/n10887_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12195_9 )
);
defparam \top/processor/sha_core/n12195_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12196_s5  (
	.I0(\top/processor/core_hash_init [194]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10888_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12196_9 )
);
defparam \top/processor/sha_core/n12196_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12197_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [193]),
	.I2(\top/processor/sha_core/n10889_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12197_9 )
);
defparam \top/processor/sha_core/n12197_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12198_s5  (
	.I0(\top/processor/core_hash_init [192]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10890_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12198_9 )
);
defparam \top/processor/sha_core/n12198_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12199_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [191]),
	.I2(\top/processor/sha_core/n10892_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12199_9 )
);
defparam \top/processor/sha_core/n12199_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12200_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [190]),
	.I2(\top/processor/sha_core/n10893_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12200_9 )
);
defparam \top/processor/sha_core/n12200_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12201_s5  (
	.I0(\top/processor/core_hash_init [189]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10894_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12201_9 )
);
defparam \top/processor/sha_core/n12201_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12202_s5  (
	.I0(\top/processor/core_hash_init [188]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10895_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12202_9 )
);
defparam \top/processor/sha_core/n12202_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12203_s5  (
	.I0(\top/processor/core_hash_init [187]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10896_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12203_9 )
);
defparam \top/processor/sha_core/n12203_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12204_s5  (
	.I0(\top/processor/core_hash_init [186]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10897_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12204_9 )
);
defparam \top/processor/sha_core/n12204_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12205_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [185]),
	.I2(\top/processor/sha_core/n10898_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12205_9 )
);
defparam \top/processor/sha_core/n12205_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12206_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [184]),
	.I2(\top/processor/sha_core/n10899_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12206_9 )
);
defparam \top/processor/sha_core/n12206_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12207_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [183]),
	.I2(\top/processor/sha_core/n10900_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12207_9 )
);
defparam \top/processor/sha_core/n12207_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12208_s5  (
	.I0(\top/processor/core_hash_init [182]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10901_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12208_9 )
);
defparam \top/processor/sha_core/n12208_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12209_s5  (
	.I0(\top/processor/core_hash_init [181]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10902_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12209_9 )
);
defparam \top/processor/sha_core/n12209_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12210_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [180]),
	.I2(\top/processor/sha_core/n10903_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12210_9 )
);
defparam \top/processor/sha_core/n12210_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12211_s5  (
	.I0(\top/processor/core_hash_init [179]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10904_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12211_9 )
);
defparam \top/processor/sha_core/n12211_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12212_s5  (
	.I0(\top/processor/core_hash_init [178]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10905_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12212_9 )
);
defparam \top/processor/sha_core/n12212_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12213_s5  (
	.I0(\top/processor/core_hash_init [177]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10906_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12213_9 )
);
defparam \top/processor/sha_core/n12213_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12214_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [176]),
	.I2(\top/processor/sha_core/n10907_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12214_9 )
);
defparam \top/processor/sha_core/n12214_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12215_s5  (
	.I0(\top/processor/core_hash_init [175]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10908_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12215_9 )
);
defparam \top/processor/sha_core/n12215_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12216_s5  (
	.I0(\top/processor/core_hash_init [174]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10909_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12216_9 )
);
defparam \top/processor/sha_core/n12216_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12217_s5  (
	.I0(\top/processor/core_hash_init [173]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10910_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12217_9 )
);
defparam \top/processor/sha_core/n12217_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12218_s5  (
	.I0(\top/processor/core_hash_init [172]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10911_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12218_9 )
);
defparam \top/processor/sha_core/n12218_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12219_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [171]),
	.I2(\top/processor/sha_core/n10912_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12219_9 )
);
defparam \top/processor/sha_core/n12219_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12220_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [170]),
	.I2(\top/processor/sha_core/n10913_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12220_9 )
);
defparam \top/processor/sha_core/n12220_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12221_s5  (
	.I0(\top/processor/core_hash_init [169]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10914_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12221_9 )
);
defparam \top/processor/sha_core/n12221_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12222_s5  (
	.I0(\top/processor/core_hash_init [168]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10915_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12222_9 )
);
defparam \top/processor/sha_core/n12222_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12223_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [167]),
	.I2(\top/processor/sha_core/n10916_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12223_9 )
);
defparam \top/processor/sha_core/n12223_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12224_s5  (
	.I0(\top/processor/core_hash_init [166]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10917_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12224_9 )
);
defparam \top/processor/sha_core/n12224_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12225_s5  (
	.I0(\top/processor/core_hash_init [165]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10918_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12225_9 )
);
defparam \top/processor/sha_core/n12225_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12226_s5  (
	.I0(\top/processor/core_hash_init [164]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10919_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12226_9 )
);
defparam \top/processor/sha_core/n12226_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12227_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [163]),
	.I2(\top/processor/sha_core/n10920_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12227_9 )
);
defparam \top/processor/sha_core/n12227_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12228_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [162]),
	.I2(\top/processor/sha_core/n10921_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12228_9 )
);
defparam \top/processor/sha_core/n12228_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12229_s5  (
	.I0(\top/processor/core_hash_init [161]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10922_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12229_9 )
);
defparam \top/processor/sha_core/n12229_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12230_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [160]),
	.I2(\top/processor/sha_core/n10923_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12230_9 )
);
defparam \top/processor/sha_core/n12230_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12231_s5  (
	.I0(\top/processor/core_hash_init [159]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10925_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12231_9 )
);
defparam \top/processor/sha_core/n12231_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12232_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [158]),
	.I2(\top/processor/sha_core/n10926_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12232_9 )
);
defparam \top/processor/sha_core/n12232_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12233_s5  (
	.I0(\top/processor/core_hash_init [157]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10927_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12233_9 )
);
defparam \top/processor/sha_core/n12233_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12234_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [156]),
	.I2(\top/processor/sha_core/n10928_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12234_9 )
);
defparam \top/processor/sha_core/n12234_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12235_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [155]),
	.I2(\top/processor/sha_core/n10929_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12235_9 )
);
defparam \top/processor/sha_core/n12235_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12236_s5  (
	.I0(\top/processor/core_hash_init [154]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10930_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12236_9 )
);
defparam \top/processor/sha_core/n12236_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12237_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [153]),
	.I2(\top/processor/sha_core/n10931_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12237_9 )
);
defparam \top/processor/sha_core/n12237_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12238_s5  (
	.I0(\top/processor/core_hash_init [152]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10932_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12238_9 )
);
defparam \top/processor/sha_core/n12238_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12239_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [151]),
	.I2(\top/processor/sha_core/n10933_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12239_9 )
);
defparam \top/processor/sha_core/n12239_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12240_s5  (
	.I0(\top/processor/core_hash_init [150]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10934_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12240_9 )
);
defparam \top/processor/sha_core/n12240_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12241_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [149]),
	.I2(\top/processor/sha_core/n10935_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12241_9 )
);
defparam \top/processor/sha_core/n12241_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12242_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [148]),
	.I2(\top/processor/sha_core/n10936_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12242_9 )
);
defparam \top/processor/sha_core/n12242_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12243_s5  (
	.I0(\top/processor/core_hash_init [147]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10937_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12243_9 )
);
defparam \top/processor/sha_core/n12243_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12244_s5  (
	.I0(\top/processor/core_hash_init [146]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10938_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12244_9 )
);
defparam \top/processor/sha_core/n12244_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12245_s5  (
	.I0(\top/processor/core_hash_init [145]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10939_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12245_9 )
);
defparam \top/processor/sha_core/n12245_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12246_s5  (
	.I0(\top/processor/core_hash_init [144]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10940_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12246_9 )
);
defparam \top/processor/sha_core/n12246_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12247_s5  (
	.I0(\top/processor/core_hash_init [143]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10941_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12247_9 )
);
defparam \top/processor/sha_core/n12247_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12248_s5  (
	.I0(\top/processor/core_hash_init [142]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10942_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12248_9 )
);
defparam \top/processor/sha_core/n12248_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12249_s5  (
	.I0(\top/processor/core_hash_init [141]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10943_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12249_9 )
);
defparam \top/processor/sha_core/n12249_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12250_s5  (
	.I0(\top/processor/core_hash_init [140]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10944_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12250_9 )
);
defparam \top/processor/sha_core/n12250_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12251_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [139]),
	.I2(\top/processor/sha_core/n10945_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12251_9 )
);
defparam \top/processor/sha_core/n12251_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12252_s5  (
	.I0(\top/processor/core_hash_init [138]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10946_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12252_9 )
);
defparam \top/processor/sha_core/n12252_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12253_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [137]),
	.I2(\top/processor/sha_core/n10947_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12253_9 )
);
defparam \top/processor/sha_core/n12253_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12254_s5  (
	.I0(\top/processor/core_hash_init [136]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10948_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12254_9 )
);
defparam \top/processor/sha_core/n12254_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12255_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [135]),
	.I2(\top/processor/sha_core/n10949_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12255_9 )
);
defparam \top/processor/sha_core/n12255_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12256_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [134]),
	.I2(\top/processor/sha_core/n10950_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12256_9 )
);
defparam \top/processor/sha_core/n12256_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12257_s5  (
	.I0(\top/processor/core_hash_init [133]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10951_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12257_9 )
);
defparam \top/processor/sha_core/n12257_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12258_s5  (
	.I0(\top/processor/core_hash_init [132]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10952_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12258_9 )
);
defparam \top/processor/sha_core/n12258_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12259_s5  (
	.I0(\top/processor/core_hash_init [131]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10953_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12259_9 )
);
defparam \top/processor/sha_core/n12259_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12260_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [130]),
	.I2(\top/processor/sha_core/n10954_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12260_9 )
);
defparam \top/processor/sha_core/n12260_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12261_s5  (
	.I0(\top/processor/core_hash_init [129]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10955_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12261_9 )
);
defparam \top/processor/sha_core/n12261_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12262_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [128]),
	.I2(\top/processor/sha_core/n10956_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12262_9 )
);
defparam \top/processor/sha_core/n12262_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12263_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [127]),
	.I2(\top/processor/sha_core/n10958_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12263_9 )
);
defparam \top/processor/sha_core/n12263_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12264_s5  (
	.I0(\top/processor/core_hash_init [126]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10959_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12264_9 )
);
defparam \top/processor/sha_core/n12264_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12265_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [125]),
	.I2(\top/processor/sha_core/n10960_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12265_9 )
);
defparam \top/processor/sha_core/n12265_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12266_s5  (
	.I0(\top/processor/core_hash_init [124]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10961_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12266_9 )
);
defparam \top/processor/sha_core/n12266_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12267_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [123]),
	.I2(\top/processor/sha_core/n10962_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12267_9 )
);
defparam \top/processor/sha_core/n12267_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12268_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [122]),
	.I2(\top/processor/sha_core/n10963_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12268_9 )
);
defparam \top/processor/sha_core/n12268_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12269_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [121]),
	.I2(\top/processor/sha_core/n10964_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12269_9 )
);
defparam \top/processor/sha_core/n12269_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12270_s5  (
	.I0(\top/processor/core_hash_init [120]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10965_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12270_9 )
);
defparam \top/processor/sha_core/n12270_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12271_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [119]),
	.I2(\top/processor/sha_core/n10966_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12271_9 )
);
defparam \top/processor/sha_core/n12271_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12272_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [118]),
	.I2(\top/processor/sha_core/n10967_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12272_9 )
);
defparam \top/processor/sha_core/n12272_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12273_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [117]),
	.I2(\top/processor/sha_core/n10968_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12273_9 )
);
defparam \top/processor/sha_core/n12273_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12274_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [116]),
	.I2(\top/processor/sha_core/n10969_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12274_9 )
);
defparam \top/processor/sha_core/n12274_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12275_s5  (
	.I0(\top/processor/core_hash_init [115]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10970_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12275_9 )
);
defparam \top/processor/sha_core/n12275_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12276_s5  (
	.I0(\top/processor/core_hash_init [114]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10971_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12276_9 )
);
defparam \top/processor/sha_core/n12276_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12277_s5  (
	.I0(\top/processor/core_hash_init [113]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10972_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12277_9 )
);
defparam \top/processor/sha_core/n12277_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12278_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [112]),
	.I2(\top/processor/sha_core/n10973_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12278_9 )
);
defparam \top/processor/sha_core/n12278_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12279_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [111]),
	.I2(\top/processor/sha_core/n10974_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12279_9 )
);
defparam \top/processor/sha_core/n12279_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12280_s5  (
	.I0(\top/processor/core_hash_init [110]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10975_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12280_9 )
);
defparam \top/processor/sha_core/n12280_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12281_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [109]),
	.I2(\top/processor/sha_core/n10976_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12281_9 )
);
defparam \top/processor/sha_core/n12281_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12282_s5  (
	.I0(\top/processor/core_hash_init [108]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10977_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12282_9 )
);
defparam \top/processor/sha_core/n12282_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12283_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [107]),
	.I2(\top/processor/sha_core/n10978_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12283_9 )
);
defparam \top/processor/sha_core/n12283_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12284_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [106]),
	.I2(\top/processor/sha_core/n10979_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12284_9 )
);
defparam \top/processor/sha_core/n12284_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12285_s5  (
	.I0(\top/processor/core_hash_init [105]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10980_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12285_9 )
);
defparam \top/processor/sha_core/n12285_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12286_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [104]),
	.I2(\top/processor/sha_core/n10981_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12286_9 )
);
defparam \top/processor/sha_core/n12286_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12287_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [103]),
	.I2(\top/processor/sha_core/n10982_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12287_9 )
);
defparam \top/processor/sha_core/n12287_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12288_s5  (
	.I0(\top/processor/core_hash_init [102]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10983_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12288_9 )
);
defparam \top/processor/sha_core/n12288_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12289_s5  (
	.I0(\top/processor/core_hash_init [101]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10984_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12289_9 )
);
defparam \top/processor/sha_core/n12289_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12290_s5  (
	.I0(\top/processor/core_hash_init [100]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10985_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12290_9 )
);
defparam \top/processor/sha_core/n12290_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12291_s5  (
	.I0(\top/processor/core_hash_init [99]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10986_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12291_9 )
);
defparam \top/processor/sha_core/n12291_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12292_s5  (
	.I0(\top/processor/core_hash_init [98]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10987_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12292_9 )
);
defparam \top/processor/sha_core/n12292_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12293_s5  (
	.I0(\top/processor/core_hash_init [97]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10988_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12293_9 )
);
defparam \top/processor/sha_core/n12293_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12294_s5  (
	.I0(\top/processor/core_hash_init [96]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10989_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12294_9 )
);
defparam \top/processor/sha_core/n12294_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12295_s5  (
	.I0(\top/processor/core_hash_init [95]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10991_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12295_9 )
);
defparam \top/processor/sha_core/n12295_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12296_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [94]),
	.I2(\top/processor/sha_core/n10992_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12296_9 )
);
defparam \top/processor/sha_core/n12296_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12297_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [93]),
	.I2(\top/processor/sha_core/n10993_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12297_9 )
);
defparam \top/processor/sha_core/n12297_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12298_s5  (
	.I0(\top/processor/core_hash_init [92]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10994_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12298_9 )
);
defparam \top/processor/sha_core/n12298_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12299_s5  (
	.I0(\top/processor/core_hash_init [91]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10995_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12299_9 )
);
defparam \top/processor/sha_core/n12299_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12300_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [90]),
	.I2(\top/processor/sha_core/n10996_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12300_9 )
);
defparam \top/processor/sha_core/n12300_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12301_s5  (
	.I0(\top/processor/core_hash_init [89]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10997_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12301_9 )
);
defparam \top/processor/sha_core/n12301_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12302_s5  (
	.I0(\top/processor/core_hash_init [88]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n10998_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12302_9 )
);
defparam \top/processor/sha_core/n12302_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12303_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [87]),
	.I2(\top/processor/sha_core/n10999_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12303_9 )
);
defparam \top/processor/sha_core/n12303_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12304_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [86]),
	.I2(\top/processor/sha_core/n11000_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12304_9 )
);
defparam \top/processor/sha_core/n12304_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12305_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [85]),
	.I2(\top/processor/sha_core/n11001_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12305_9 )
);
defparam \top/processor/sha_core/n12305_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12306_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [84]),
	.I2(\top/processor/sha_core/n11002_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12306_9 )
);
defparam \top/processor/sha_core/n12306_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12307_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [83]),
	.I2(\top/processor/sha_core/n11003_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12307_9 )
);
defparam \top/processor/sha_core/n12307_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12308_s5  (
	.I0(\top/processor/core_hash_init [82]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11004_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12308_9 )
);
defparam \top/processor/sha_core/n12308_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12309_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [81]),
	.I2(\top/processor/sha_core/n11005_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12309_9 )
);
defparam \top/processor/sha_core/n12309_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12310_s5  (
	.I0(\top/processor/core_hash_init [80]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11006_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12310_9 )
);
defparam \top/processor/sha_core/n12310_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12311_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [79]),
	.I2(\top/processor/sha_core/n11007_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12311_9 )
);
defparam \top/processor/sha_core/n12311_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12312_s5  (
	.I0(\top/processor/core_hash_init [78]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11008_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12312_9 )
);
defparam \top/processor/sha_core/n12312_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12313_s5  (
	.I0(\top/processor/core_hash_init [77]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11009_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12313_9 )
);
defparam \top/processor/sha_core/n12313_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12314_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [76]),
	.I2(\top/processor/sha_core/n11010_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12314_9 )
);
defparam \top/processor/sha_core/n12314_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12315_s5  (
	.I0(\top/processor/core_hash_init [75]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11011_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12315_9 )
);
defparam \top/processor/sha_core/n12315_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12316_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [74]),
	.I2(\top/processor/sha_core/n11012_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12316_9 )
);
defparam \top/processor/sha_core/n12316_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12317_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [73]),
	.I2(\top/processor/sha_core/n11013_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12317_9 )
);
defparam \top/processor/sha_core/n12317_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12318_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [72]),
	.I2(\top/processor/sha_core/n11014_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12318_9 )
);
defparam \top/processor/sha_core/n12318_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12319_s5  (
	.I0(\top/processor/core_hash_init [71]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11015_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12319_9 )
);
defparam \top/processor/sha_core/n12319_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12320_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [70]),
	.I2(\top/processor/sha_core/n11016_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12320_9 )
);
defparam \top/processor/sha_core/n12320_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12321_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [69]),
	.I2(\top/processor/sha_core/n11017_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12321_9 )
);
defparam \top/processor/sha_core/n12321_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12322_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [68]),
	.I2(\top/processor/sha_core/n11018_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12322_9 )
);
defparam \top/processor/sha_core/n12322_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12323_s5  (
	.I0(\top/processor/core_hash_init [67]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11019_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12323_9 )
);
defparam \top/processor/sha_core/n12323_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12324_s5  (
	.I0(\top/processor/core_hash_init [66]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11020_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12324_9 )
);
defparam \top/processor/sha_core/n12324_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12325_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [65]),
	.I2(\top/processor/sha_core/n11021_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12325_9 )
);
defparam \top/processor/sha_core/n12325_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12326_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [64]),
	.I2(\top/processor/sha_core/n11022_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12326_9 )
);
defparam \top/processor/sha_core/n12326_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12327_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [63]),
	.I2(\top/processor/sha_core/n11024_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12327_9 )
);
defparam \top/processor/sha_core/n12327_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12328_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [62]),
	.I2(\top/processor/sha_core/n11025_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12328_9 )
);
defparam \top/processor/sha_core/n12328_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12329_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [61]),
	.I2(\top/processor/sha_core/n11026_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12329_9 )
);
defparam \top/processor/sha_core/n12329_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12330_s5  (
	.I0(\top/processor/core_hash_init [60]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11027_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12330_9 )
);
defparam \top/processor/sha_core/n12330_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12331_s5  (
	.I0(\top/processor/core_hash_init [59]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11028_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12331_9 )
);
defparam \top/processor/sha_core/n12331_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12332_s5  (
	.I0(\top/processor/core_hash_init [58]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11029_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12332_9 )
);
defparam \top/processor/sha_core/n12332_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12333_s5  (
	.I0(\top/processor/core_hash_init [57]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11030_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12333_9 )
);
defparam \top/processor/sha_core/n12333_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12334_s5  (
	.I0(\top/processor/core_hash_init [56]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11031_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12334_9 )
);
defparam \top/processor/sha_core/n12334_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12335_s5  (
	.I0(\top/processor/core_hash_init [55]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11032_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12335_9 )
);
defparam \top/processor/sha_core/n12335_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12336_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [54]),
	.I2(\top/processor/sha_core/n11033_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12336_9 )
);
defparam \top/processor/sha_core/n12336_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12337_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [53]),
	.I2(\top/processor/sha_core/n11034_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12337_9 )
);
defparam \top/processor/sha_core/n12337_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12338_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [52]),
	.I2(\top/processor/sha_core/n11035_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12338_9 )
);
defparam \top/processor/sha_core/n12338_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12339_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [51]),
	.I2(\top/processor/sha_core/n11036_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12339_9 )
);
defparam \top/processor/sha_core/n12339_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12340_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [50]),
	.I2(\top/processor/sha_core/n11037_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12340_9 )
);
defparam \top/processor/sha_core/n12340_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12341_s5  (
	.I0(\top/processor/core_hash_init [49]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11038_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12341_9 )
);
defparam \top/processor/sha_core/n12341_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12342_s5  (
	.I0(\top/processor/core_hash_init [48]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11039_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12342_9 )
);
defparam \top/processor/sha_core/n12342_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12343_s5  (
	.I0(\top/processor/core_hash_init [47]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11040_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12343_9 )
);
defparam \top/processor/sha_core/n12343_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12344_s5  (
	.I0(\top/processor/core_hash_init [46]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11041_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12344_9 )
);
defparam \top/processor/sha_core/n12344_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12345_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [45]),
	.I2(\top/processor/sha_core/n11042_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12345_9 )
);
defparam \top/processor/sha_core/n12345_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12346_s5  (
	.I0(\top/processor/core_hash_init [44]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11043_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12346_9 )
);
defparam \top/processor/sha_core/n12346_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12347_s5  (
	.I0(\top/processor/core_hash_init [43]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11044_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12347_9 )
);
defparam \top/processor/sha_core/n12347_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12348_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [42]),
	.I2(\top/processor/sha_core/n11045_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12348_9 )
);
defparam \top/processor/sha_core/n12348_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12349_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [41]),
	.I2(\top/processor/sha_core/n11046_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12349_9 )
);
defparam \top/processor/sha_core/n12349_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12350_s5  (
	.I0(\top/processor/core_hash_init [40]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11047_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12350_9 )
);
defparam \top/processor/sha_core/n12350_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12351_s5  (
	.I0(\top/processor/core_hash_init [39]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11048_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12351_9 )
);
defparam \top/processor/sha_core/n12351_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12352_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [38]),
	.I2(\top/processor/sha_core/n11049_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12352_9 )
);
defparam \top/processor/sha_core/n12352_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12353_s5  (
	.I0(\top/processor/core_hash_init [37]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11050_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12353_9 )
);
defparam \top/processor/sha_core/n12353_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12354_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [36]),
	.I2(\top/processor/sha_core/n11051_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12354_9 )
);
defparam \top/processor/sha_core/n12354_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12355_s5  (
	.I0(\top/processor/core_hash_init [35]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11052_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12355_9 )
);
defparam \top/processor/sha_core/n12355_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12356_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [34]),
	.I2(\top/processor/sha_core/n11053_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12356_9 )
);
defparam \top/processor/sha_core/n12356_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12357_s5  (
	.I0(\top/processor/core_hash_init [33]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11054_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12357_9 )
);
defparam \top/processor/sha_core/n12357_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12358_s5  (
	.I0(\top/processor/core_hash_init [32]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11055_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12358_9 )
);
defparam \top/processor/sha_core/n12358_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12359_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [31]),
	.I2(\top/processor/sha_core/n11057_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12359_9 )
);
defparam \top/processor/sha_core/n12359_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12360_s5  (
	.I0(\top/processor/core_hash_init [30]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11058_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12360_9 )
);
defparam \top/processor/sha_core/n12360_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12361_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [29]),
	.I2(\top/processor/sha_core/n11059_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12361_9 )
);
defparam \top/processor/sha_core/n12361_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12362_s5  (
	.I0(\top/processor/core_hash_init [28]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11060_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12362_9 )
);
defparam \top/processor/sha_core/n12362_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12363_s5  (
	.I0(\top/processor/core_hash_init [27]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11061_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12363_9 )
);
defparam \top/processor/sha_core/n12363_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12364_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [26]),
	.I2(\top/processor/sha_core/n11062_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12364_9 )
);
defparam \top/processor/sha_core/n12364_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12365_s5  (
	.I0(\top/processor/core_hash_init [25]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11063_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12365_9 )
);
defparam \top/processor/sha_core/n12365_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12366_s5  (
	.I0(\top/processor/core_hash_init [24]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11064_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12366_9 )
);
defparam \top/processor/sha_core/n12366_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12367_s5  (
	.I0(\top/processor/core_hash_init [23]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11065_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12367_9 )
);
defparam \top/processor/sha_core/n12367_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12368_s5  (
	.I0(\top/processor/core_hash_init [22]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11066_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12368_9 )
);
defparam \top/processor/sha_core/n12368_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12369_s5  (
	.I0(\top/processor/core_hash_init [21]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11067_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12369_9 )
);
defparam \top/processor/sha_core/n12369_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12370_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [20]),
	.I2(\top/processor/sha_core/n11068_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12370_9 )
);
defparam \top/processor/sha_core/n12370_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12371_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [19]),
	.I2(\top/processor/sha_core/n11069_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12371_9 )
);
defparam \top/processor/sha_core/n12371_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12372_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [18]),
	.I2(\top/processor/sha_core/n11070_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12372_9 )
);
defparam \top/processor/sha_core/n12372_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12373_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [17]),
	.I2(\top/processor/sha_core/n11071_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12373_9 )
);
defparam \top/processor/sha_core/n12373_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12374_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [16]),
	.I2(\top/processor/sha_core/n11072_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12374_9 )
);
defparam \top/processor/sha_core/n12374_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12375_s5  (
	.I0(\top/processor/core_hash_init [15]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11073_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12375_9 )
);
defparam \top/processor/sha_core/n12375_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12376_s5  (
	.I0(\top/processor/core_hash_init [14]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11074_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12376_9 )
);
defparam \top/processor/sha_core/n12376_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12377_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [13]),
	.I2(\top/processor/sha_core/n11075_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12377_9 )
);
defparam \top/processor/sha_core/n12377_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12378_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [12]),
	.I2(\top/processor/sha_core/n11076_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12378_9 )
);
defparam \top/processor/sha_core/n12378_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12379_s5  (
	.I0(\top/processor/core_hash_init [11]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11077_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12379_9 )
);
defparam \top/processor/sha_core/n12379_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12380_s5  (
	.I0(\top/processor/core_hash_init [10]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11078_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12380_9 )
);
defparam \top/processor/sha_core/n12380_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12381_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [9]),
	.I2(\top/processor/sha_core/n11079_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12381_9 )
);
defparam \top/processor/sha_core/n12381_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12382_s5  (
	.I0(\top/processor/core_hash_init [8]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11080_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12382_9 )
);
defparam \top/processor/sha_core/n12382_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12383_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [7]),
	.I2(\top/processor/sha_core/n11081_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12383_9 )
);
defparam \top/processor/sha_core/n12383_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12384_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [6]),
	.I2(\top/processor/sha_core/n11082_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12384_9 )
);
defparam \top/processor/sha_core/n12384_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12385_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [5]),
	.I2(\top/processor/sha_core/n11083_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12385_9 )
);
defparam \top/processor/sha_core/n12385_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12386_s5  (
	.I0(\top/processor/core_hash_init [4]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11084_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12386_9 )
);
defparam \top/processor/sha_core/n12386_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12387_s5  (
	.I0(\top/processor/core_hash_init [3]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11085_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12387_9 )
);
defparam \top/processor/sha_core/n12387_s5 .INIT=16'hF0BB;
LUT4 \top/processor/sha_core/n12388_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [2]),
	.I2(\top/processor/sha_core/n11086_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12388_9 )
);
defparam \top/processor/sha_core/n12388_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12389_s5  (
	.I0(\top/processor/core_use_init ),
	.I1(\top/processor/core_hash_init [1]),
	.I2(\top/processor/sha_core/n11087_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12389_9 )
);
defparam \top/processor/sha_core/n12389_s5 .INIT=16'hF088;
LUT4 \top/processor/sha_core/n12390_s5  (
	.I0(\top/processor/core_hash_init [0]),
	.I1(\top/processor/core_use_init ),
	.I2(\top/processor/sha_core/n11088_1 ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12390_9 )
);
defparam \top/processor/sha_core/n12390_s5 .INIT=16'hF0BB;
LUT2 \top/processor/sha_core/n11613_s4  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11613_8 )
);
defparam \top/processor/sha_core/n11613_s4 .INIT=4'h8;
LUT4 \top/processor/sha_core/t_6_s3  (
	.I0(\top/processor/sha_core/t [6]),
	.I1(\top/processor/sha_core/msg_idx [6]),
	.I2(\top/processor/sha_core/state [0]),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/t_6_8 )
);
defparam \top/processor/sha_core/t_6_s3 .INIT=16'h05C0;
LUT4 \top/processor/sha_core/msg_idx_6_s3  (
	.I0(\top/processor/core_start ),
	.I1(\top/processor/sha_core/msg_idx [6]),
	.I2(\top/processor/sha_core/state [1]),
	.I3(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/msg_idx_6_7 )
);
defparam \top/processor/sha_core/msg_idx_6_s3 .INIT=16'h030A;
LUT4 \top/processor/sha_core/h0_31_s3  (
	.I0(\top/processor/sha_core/t [6]),
	.I1(\top/processor/core_start ),
	.I2(\top/processor/sha_core/state [0]),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/h0_31_8 )
);
defparam \top/processor/sha_core/h0_31_s3 .INIT=16'h0A0C;
LUT2 \top/processor/sha_core/w[2]_31_s4  (
	.I0(\top/processor/sha_core/w[2]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[2]_31_8 )
);
defparam \top/processor/sha_core/w[2]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[3]_31_s4  (
	.I0(\top/processor/sha_core/w[3]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[3]_31_8 )
);
defparam \top/processor/sha_core/w[3]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[4]_31_s4  (
	.I0(\top/processor/sha_core/w[4]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[4]_31_8 )
);
defparam \top/processor/sha_core/w[4]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[5]_31_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[5]_31_8 )
);
defparam \top/processor/sha_core/w[5]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[6]_31_s4  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[6]_31_8 )
);
defparam \top/processor/sha_core/w[6]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[7]_31_s4  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[7]_31_8 )
);
defparam \top/processor/sha_core/w[7]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[8]_31_s4  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[8]_31_8 )
);
defparam \top/processor/sha_core/w[8]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[9]_31_s4  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[9]_31_8 )
);
defparam \top/processor/sha_core/w[9]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[10]_31_s4  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[10]_31_8 )
);
defparam \top/processor/sha_core/w[10]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[11]_31_s4  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[11]_31_8 )
);
defparam \top/processor/sha_core/w[11]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[12]_31_s4  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[12]_31_8 )
);
defparam \top/processor/sha_core/w[12]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[13]_31_s4  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[13]_31_8 )
);
defparam \top/processor/sha_core/w[13]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[14]_31_s4  (
	.I0(\top/processor/sha_core/w[14]_31_9 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[14]_31_8 )
);
defparam \top/processor/sha_core/w[14]_31_s4 .INIT=4'h8;
LUT2 \top/processor/sha_core/w[15]_31_s4  (
	.I0(\top/processor/sha_core/w[15]_31_11 ),
	.I1(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[15]_31_8 )
);
defparam \top/processor/sha_core/w[15]_31_s4 .INIT=4'h8;
LUT4 \top/processor/sha_core/w[16]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[16]_31_8 )
);
defparam \top/processor/sha_core/w[16]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[17]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[17]_31_8 )
);
defparam \top/processor/sha_core/w[17]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[18]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[18]_31_9 ),
	.F(\top/processor/sha_core/w[18]_31_8 )
);
defparam \top/processor/sha_core/w[18]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[19]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[19]_31_9 ),
	.F(\top/processor/sha_core/w[19]_31_8 )
);
defparam \top/processor/sha_core/w[19]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[20]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[20]_31_9 ),
	.F(\top/processor/sha_core/w[20]_31_8 )
);
defparam \top/processor/sha_core/w[20]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[21]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[21]_31_9 ),
	.F(\top/processor/sha_core/w[21]_31_8 )
);
defparam \top/processor/sha_core/w[21]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[22]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[22]_31_9 ),
	.F(\top/processor/sha_core/w[22]_31_8 )
);
defparam \top/processor/sha_core/w[22]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[23]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[23]_31_11 ),
	.F(\top/processor/sha_core/w[23]_31_8 )
);
defparam \top/processor/sha_core/w[23]_31_s4 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[24]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[24]_31_8 )
);
defparam \top/processor/sha_core/w[24]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[25]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[25]_31_8 )
);
defparam \top/processor/sha_core/w[25]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[26]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[18]_31_9 ),
	.F(\top/processor/sha_core/w[26]_31_8 )
);
defparam \top/processor/sha_core/w[26]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[27]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[19]_31_9 ),
	.F(\top/processor/sha_core/w[27]_31_8 )
);
defparam \top/processor/sha_core/w[27]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[28]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[20]_31_9 ),
	.F(\top/processor/sha_core/w[28]_31_8 )
);
defparam \top/processor/sha_core/w[28]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[29]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[21]_31_9 ),
	.F(\top/processor/sha_core/w[29]_31_8 )
);
defparam \top/processor/sha_core/w[29]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[30]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.I3(\top/processor/sha_core/w[22]_31_9 ),
	.F(\top/processor/sha_core/w[30]_31_8 )
);
defparam \top/processor/sha_core/w[30]_31_s4 .INIT=16'h4000;
LUT3 \top/processor/sha_core/w[31]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/w[31]_31_11 ),
	.I2(\top/processor/sha_core/w[2]_31_12 ),
	.F(\top/processor/sha_core/w[31]_31_8 )
);
defparam \top/processor/sha_core/w[31]_31_s4 .INIT=8'h80;
LUT4 \top/processor/sha_core/w[48]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[48]_31_8 )
);
defparam \top/processor/sha_core/w[48]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[49]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[49]_31_8 )
);
defparam \top/processor/sha_core/w[49]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[50]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[18]_31_9 ),
	.F(\top/processor/sha_core/w[50]_31_8 )
);
defparam \top/processor/sha_core/w[50]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[51]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[19]_31_9 ),
	.F(\top/processor/sha_core/w[51]_31_8 )
);
defparam \top/processor/sha_core/w[51]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[52]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[20]_31_9 ),
	.F(\top/processor/sha_core/w[52]_31_8 )
);
defparam \top/processor/sha_core/w[52]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[53]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[21]_31_9 ),
	.F(\top/processor/sha_core/w[53]_31_8 )
);
defparam \top/processor/sha_core/w[53]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[54]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[22]_31_9 ),
	.F(\top/processor/sha_core/w[54]_31_8 )
);
defparam \top/processor/sha_core/w[54]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[55]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[23]_31_11 ),
	.F(\top/processor/sha_core/w[55]_31_8 )
);
defparam \top/processor/sha_core/w[55]_31_s4 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[56]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[56]_31_8 )
);
defparam \top/processor/sha_core/w[56]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[57]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[57]_31_8 )
);
defparam \top/processor/sha_core/w[57]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[58]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[18]_31_9 ),
	.F(\top/processor/sha_core/w[58]_31_8 )
);
defparam \top/processor/sha_core/w[58]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[59]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[19]_31_9 ),
	.F(\top/processor/sha_core/w[59]_31_8 )
);
defparam \top/processor/sha_core/w[59]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[60]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[20]_31_9 ),
	.F(\top/processor/sha_core/w[60]_31_8 )
);
defparam \top/processor/sha_core/w[60]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[61]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[21]_31_9 ),
	.F(\top/processor/sha_core/w[61]_31_8 )
);
defparam \top/processor/sha_core/w[61]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[62]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/w[22]_31_9 ),
	.F(\top/processor/sha_core/w[62]_31_8 )
);
defparam \top/processor/sha_core/w[62]_31_s4 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[63]_31_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/w[31]_31_11 ),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[63]_31_8 )
);
defparam \top/processor/sha_core/w[63]_31_s4 .INIT=16'h8000;
LUT2 \top/processor/sha_core/h_31_s4  (
	.I0(rst),
	.I1(\top/processor/sha_core/t_6_8 ),
	.F(\top/processor/sha_core/h_31_8 )
);
defparam \top/processor/sha_core/h_31_s4 .INIT=4'h4;
LUT2 \top/processor/sha_core/n3453_s3  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.F(\top/processor/sha_core/n3453_7 )
);
defparam \top/processor/sha_core/n3453_s3 .INIT=4'h6;
LUT3 \top/processor/sha_core/n3452_s3  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.F(\top/processor/sha_core/n3452_7 )
);
defparam \top/processor/sha_core/n3452_s3 .INIT=8'h78;
LUT3 \top/processor/sha_core/n327_s189  (
	.I0(\top/processor/sha_core/n327_221 ),
	.I1(\top/processor/sha_core/n327_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n327_225 )
);
defparam \top/processor/sha_core/n327_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n328_s189  (
	.I0(\top/processor/sha_core/n328_221 ),
	.I1(\top/processor/sha_core/n328_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n328_225 )
);
defparam \top/processor/sha_core/n328_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n329_s189  (
	.I0(\top/processor/sha_core/n329_221 ),
	.I1(\top/processor/sha_core/n329_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n329_225 )
);
defparam \top/processor/sha_core/n329_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n330_s189  (
	.I0(\top/processor/sha_core/n330_221 ),
	.I1(\top/processor/sha_core/n330_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n330_225 )
);
defparam \top/processor/sha_core/n330_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n331_s189  (
	.I0(\top/processor/sha_core/n331_221 ),
	.I1(\top/processor/sha_core/n331_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n331_225 )
);
defparam \top/processor/sha_core/n331_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n332_s189  (
	.I0(\top/processor/sha_core/n332_221 ),
	.I1(\top/processor/sha_core/n332_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n332_225 )
);
defparam \top/processor/sha_core/n332_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n333_s189  (
	.I0(\top/processor/sha_core/n333_221 ),
	.I1(\top/processor/sha_core/n333_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n333_225 )
);
defparam \top/processor/sha_core/n333_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n334_s189  (
	.I0(\top/processor/sha_core/n334_221 ),
	.I1(\top/processor/sha_core/n334_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n334_225 )
);
defparam \top/processor/sha_core/n334_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n335_s189  (
	.I0(\top/processor/sha_core/n335_221 ),
	.I1(\top/processor/sha_core/n335_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n335_225 )
);
defparam \top/processor/sha_core/n335_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n336_s189  (
	.I0(\top/processor/sha_core/n336_221 ),
	.I1(\top/processor/sha_core/n336_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n336_225 )
);
defparam \top/processor/sha_core/n336_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n337_s189  (
	.I0(\top/processor/sha_core/n337_221 ),
	.I1(\top/processor/sha_core/n337_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n337_225 )
);
defparam \top/processor/sha_core/n337_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n338_s189  (
	.I0(\top/processor/sha_core/n338_221 ),
	.I1(\top/processor/sha_core/n338_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n338_225 )
);
defparam \top/processor/sha_core/n338_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n339_s189  (
	.I0(\top/processor/sha_core/n339_221 ),
	.I1(\top/processor/sha_core/n339_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n339_225 )
);
defparam \top/processor/sha_core/n339_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n340_s189  (
	.I0(\top/processor/sha_core/n340_221 ),
	.I1(\top/processor/sha_core/n340_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n340_225 )
);
defparam \top/processor/sha_core/n340_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n341_s189  (
	.I0(\top/processor/sha_core/n341_221 ),
	.I1(\top/processor/sha_core/n341_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n341_225 )
);
defparam \top/processor/sha_core/n341_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n342_s189  (
	.I0(\top/processor/sha_core/n342_221 ),
	.I1(\top/processor/sha_core/n342_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n342_225 )
);
defparam \top/processor/sha_core/n342_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n343_s189  (
	.I0(\top/processor/sha_core/n343_221 ),
	.I1(\top/processor/sha_core/n343_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n343_225 )
);
defparam \top/processor/sha_core/n343_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n344_s189  (
	.I0(\top/processor/sha_core/n344_221 ),
	.I1(\top/processor/sha_core/n344_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n344_225 )
);
defparam \top/processor/sha_core/n344_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n345_s189  (
	.I0(\top/processor/sha_core/n345_221 ),
	.I1(\top/processor/sha_core/n345_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n345_225 )
);
defparam \top/processor/sha_core/n345_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n346_s189  (
	.I0(\top/processor/sha_core/n346_221 ),
	.I1(\top/processor/sha_core/n346_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n346_225 )
);
defparam \top/processor/sha_core/n346_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n347_s189  (
	.I0(\top/processor/sha_core/n347_221 ),
	.I1(\top/processor/sha_core/n347_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n347_225 )
);
defparam \top/processor/sha_core/n347_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n348_s189  (
	.I0(\top/processor/sha_core/n348_221 ),
	.I1(\top/processor/sha_core/n348_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n348_225 )
);
defparam \top/processor/sha_core/n348_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n349_s189  (
	.I0(\top/processor/sha_core/n349_221 ),
	.I1(\top/processor/sha_core/n349_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n349_225 )
);
defparam \top/processor/sha_core/n349_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n350_s189  (
	.I0(\top/processor/sha_core/n350_221 ),
	.I1(\top/processor/sha_core/n350_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n350_225 )
);
defparam \top/processor/sha_core/n350_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n351_s189  (
	.I0(\top/processor/sha_core/n351_221 ),
	.I1(\top/processor/sha_core/n351_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n351_225 )
);
defparam \top/processor/sha_core/n351_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n352_s189  (
	.I0(\top/processor/sha_core/n352_221 ),
	.I1(\top/processor/sha_core/n352_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n352_225 )
);
defparam \top/processor/sha_core/n352_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n353_s189  (
	.I0(\top/processor/sha_core/n353_221 ),
	.I1(\top/processor/sha_core/n353_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n353_225 )
);
defparam \top/processor/sha_core/n353_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n354_s189  (
	.I0(\top/processor/sha_core/n354_221 ),
	.I1(\top/processor/sha_core/n354_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n354_225 )
);
defparam \top/processor/sha_core/n354_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n355_s189  (
	.I0(\top/processor/sha_core/n355_221 ),
	.I1(\top/processor/sha_core/n355_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n355_225 )
);
defparam \top/processor/sha_core/n355_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n356_s189  (
	.I0(\top/processor/sha_core/n356_221 ),
	.I1(\top/processor/sha_core/n356_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n356_225 )
);
defparam \top/processor/sha_core/n356_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n357_s189  (
	.I0(\top/processor/sha_core/n357_221 ),
	.I1(\top/processor/sha_core/n357_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n357_225 )
);
defparam \top/processor/sha_core/n357_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n358_s189  (
	.I0(\top/processor/sha_core/n358_221 ),
	.I1(\top/processor/sha_core/n358_223 ),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n358_225 )
);
defparam \top/processor/sha_core/n358_s189 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n3607_s170  (
	.I0(\top/processor/sha_core/n3705_135 ),
	.I1(\top/processor/sha_core/n3705_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3607_187 )
);
defparam \top/processor/sha_core/n3607_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3607_s171  (
	.I0(\top/processor/sha_core/n3705_139 ),
	.I1(\top/processor/sha_core/n3705_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3607_189 )
);
defparam \top/processor/sha_core/n3607_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3607_s172  (
	.I0(\top/processor/sha_core/n3705_143 ),
	.I1(\top/processor/sha_core/n3705_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3607_191 )
);
defparam \top/processor/sha_core/n3607_s172 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3607_s173  (
	.I0(\top/processor/sha_core/n3705_147 ),
	.I1(\top/processor/sha_core/n3705_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3607_193 )
);
defparam \top/processor/sha_core/n3607_s173 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3608_s168  (
	.I0(\top/processor/sha_core/n3706_135 ),
	.I1(\top/processor/sha_core/n3706_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3608_187 )
);
defparam \top/processor/sha_core/n3608_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3608_s169  (
	.I0(\top/processor/sha_core/n3706_139 ),
	.I1(\top/processor/sha_core/n3706_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3608_189 )
);
defparam \top/processor/sha_core/n3608_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3608_s170  (
	.I0(\top/processor/sha_core/n3706_143 ),
	.I1(\top/processor/sha_core/n3706_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3608_191 )
);
defparam \top/processor/sha_core/n3608_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3608_s171  (
	.I0(\top/processor/sha_core/n3706_147 ),
	.I1(\top/processor/sha_core/n3706_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3608_193 )
);
defparam \top/processor/sha_core/n3608_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3609_s168  (
	.I0(\top/processor/sha_core/n3707_135 ),
	.I1(\top/processor/sha_core/n3707_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3609_187 )
);
defparam \top/processor/sha_core/n3609_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3609_s169  (
	.I0(\top/processor/sha_core/n3707_139 ),
	.I1(\top/processor/sha_core/n3707_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3609_189 )
);
defparam \top/processor/sha_core/n3609_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3609_s170  (
	.I0(\top/processor/sha_core/n3707_143 ),
	.I1(\top/processor/sha_core/n3707_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3609_191 )
);
defparam \top/processor/sha_core/n3609_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3609_s171  (
	.I0(\top/processor/sha_core/n3707_147 ),
	.I1(\top/processor/sha_core/n3707_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3609_193 )
);
defparam \top/processor/sha_core/n3609_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3610_s168  (
	.I0(\top/processor/sha_core/n3708_135 ),
	.I1(\top/processor/sha_core/n3708_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3610_187 )
);
defparam \top/processor/sha_core/n3610_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3610_s169  (
	.I0(\top/processor/sha_core/n3708_139 ),
	.I1(\top/processor/sha_core/n3708_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3610_189 )
);
defparam \top/processor/sha_core/n3610_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3610_s170  (
	.I0(\top/processor/sha_core/n3708_143 ),
	.I1(\top/processor/sha_core/n3708_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3610_191 )
);
defparam \top/processor/sha_core/n3610_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3610_s171  (
	.I0(\top/processor/sha_core/n3708_147 ),
	.I1(\top/processor/sha_core/n3708_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3610_193 )
);
defparam \top/processor/sha_core/n3610_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3611_s168  (
	.I0(\top/processor/sha_core/n3709_135 ),
	.I1(\top/processor/sha_core/n3709_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3611_187 )
);
defparam \top/processor/sha_core/n3611_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3611_s169  (
	.I0(\top/processor/sha_core/n3709_139 ),
	.I1(\top/processor/sha_core/n3709_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3611_189 )
);
defparam \top/processor/sha_core/n3611_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3611_s170  (
	.I0(\top/processor/sha_core/n3709_143 ),
	.I1(\top/processor/sha_core/n3709_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3611_191 )
);
defparam \top/processor/sha_core/n3611_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3611_s171  (
	.I0(\top/processor/sha_core/n3709_147 ),
	.I1(\top/processor/sha_core/n3709_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3611_193 )
);
defparam \top/processor/sha_core/n3611_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3612_s168  (
	.I0(\top/processor/sha_core/n3710_135 ),
	.I1(\top/processor/sha_core/n3710_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3612_187 )
);
defparam \top/processor/sha_core/n3612_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3612_s169  (
	.I0(\top/processor/sha_core/n3710_139 ),
	.I1(\top/processor/sha_core/n3710_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3612_189 )
);
defparam \top/processor/sha_core/n3612_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3612_s170  (
	.I0(\top/processor/sha_core/n3710_143 ),
	.I1(\top/processor/sha_core/n3710_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3612_191 )
);
defparam \top/processor/sha_core/n3612_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3612_s171  (
	.I0(\top/processor/sha_core/n3710_147 ),
	.I1(\top/processor/sha_core/n3710_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3612_193 )
);
defparam \top/processor/sha_core/n3612_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3613_s168  (
	.I0(\top/processor/sha_core/n3711_135 ),
	.I1(\top/processor/sha_core/n3711_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3613_187 )
);
defparam \top/processor/sha_core/n3613_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3613_s169  (
	.I0(\top/processor/sha_core/n3711_139 ),
	.I1(\top/processor/sha_core/n3711_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3613_189 )
);
defparam \top/processor/sha_core/n3613_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3613_s170  (
	.I0(\top/processor/sha_core/n3711_143 ),
	.I1(\top/processor/sha_core/n3711_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3613_191 )
);
defparam \top/processor/sha_core/n3613_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3613_s171  (
	.I0(\top/processor/sha_core/n3711_147 ),
	.I1(\top/processor/sha_core/n3711_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3613_193 )
);
defparam \top/processor/sha_core/n3613_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3614_s168  (
	.I0(\top/processor/sha_core/n3712_135 ),
	.I1(\top/processor/sha_core/n3712_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3614_187 )
);
defparam \top/processor/sha_core/n3614_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3614_s169  (
	.I0(\top/processor/sha_core/n3712_139 ),
	.I1(\top/processor/sha_core/n3712_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3614_189 )
);
defparam \top/processor/sha_core/n3614_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3614_s170  (
	.I0(\top/processor/sha_core/n3712_143 ),
	.I1(\top/processor/sha_core/n3712_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3614_191 )
);
defparam \top/processor/sha_core/n3614_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3614_s171  (
	.I0(\top/processor/sha_core/n3712_147 ),
	.I1(\top/processor/sha_core/n3712_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3614_193 )
);
defparam \top/processor/sha_core/n3614_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3615_s168  (
	.I0(\top/processor/sha_core/n3713_135 ),
	.I1(\top/processor/sha_core/n3713_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3615_187 )
);
defparam \top/processor/sha_core/n3615_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3615_s169  (
	.I0(\top/processor/sha_core/n3713_139 ),
	.I1(\top/processor/sha_core/n3713_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3615_189 )
);
defparam \top/processor/sha_core/n3615_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3615_s170  (
	.I0(\top/processor/sha_core/n3713_143 ),
	.I1(\top/processor/sha_core/n3713_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3615_191 )
);
defparam \top/processor/sha_core/n3615_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3615_s171  (
	.I0(\top/processor/sha_core/n3713_147 ),
	.I1(\top/processor/sha_core/n3713_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3615_193 )
);
defparam \top/processor/sha_core/n3615_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3616_s168  (
	.I0(\top/processor/sha_core/n3714_135 ),
	.I1(\top/processor/sha_core/n3714_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3616_187 )
);
defparam \top/processor/sha_core/n3616_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3616_s169  (
	.I0(\top/processor/sha_core/n3714_139 ),
	.I1(\top/processor/sha_core/n3714_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3616_189 )
);
defparam \top/processor/sha_core/n3616_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3616_s170  (
	.I0(\top/processor/sha_core/n3714_143 ),
	.I1(\top/processor/sha_core/n3714_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3616_191 )
);
defparam \top/processor/sha_core/n3616_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3616_s171  (
	.I0(\top/processor/sha_core/n3714_147 ),
	.I1(\top/processor/sha_core/n3714_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3616_193 )
);
defparam \top/processor/sha_core/n3616_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3617_s168  (
	.I0(\top/processor/sha_core/n3715_135 ),
	.I1(\top/processor/sha_core/n3715_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3617_187 )
);
defparam \top/processor/sha_core/n3617_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3617_s169  (
	.I0(\top/processor/sha_core/n3715_139 ),
	.I1(\top/processor/sha_core/n3715_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3617_189 )
);
defparam \top/processor/sha_core/n3617_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3617_s170  (
	.I0(\top/processor/sha_core/n3715_143 ),
	.I1(\top/processor/sha_core/n3715_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3617_191 )
);
defparam \top/processor/sha_core/n3617_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3617_s171  (
	.I0(\top/processor/sha_core/n3715_147 ),
	.I1(\top/processor/sha_core/n3715_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3617_193 )
);
defparam \top/processor/sha_core/n3617_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3618_s168  (
	.I0(\top/processor/sha_core/n3716_135 ),
	.I1(\top/processor/sha_core/n3716_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3618_187 )
);
defparam \top/processor/sha_core/n3618_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3618_s169  (
	.I0(\top/processor/sha_core/n3716_139 ),
	.I1(\top/processor/sha_core/n3716_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3618_189 )
);
defparam \top/processor/sha_core/n3618_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3618_s170  (
	.I0(\top/processor/sha_core/n3716_143 ),
	.I1(\top/processor/sha_core/n3716_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3618_191 )
);
defparam \top/processor/sha_core/n3618_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3618_s171  (
	.I0(\top/processor/sha_core/n3716_147 ),
	.I1(\top/processor/sha_core/n3716_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3618_193 )
);
defparam \top/processor/sha_core/n3618_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3619_s168  (
	.I0(\top/processor/sha_core/n3717_135 ),
	.I1(\top/processor/sha_core/n3717_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3619_187 )
);
defparam \top/processor/sha_core/n3619_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3619_s169  (
	.I0(\top/processor/sha_core/n3717_139 ),
	.I1(\top/processor/sha_core/n3717_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3619_189 )
);
defparam \top/processor/sha_core/n3619_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3619_s170  (
	.I0(\top/processor/sha_core/n3717_143 ),
	.I1(\top/processor/sha_core/n3717_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3619_191 )
);
defparam \top/processor/sha_core/n3619_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3619_s171  (
	.I0(\top/processor/sha_core/n3717_147 ),
	.I1(\top/processor/sha_core/n3717_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3619_193 )
);
defparam \top/processor/sha_core/n3619_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3620_s168  (
	.I0(\top/processor/sha_core/n3718_135 ),
	.I1(\top/processor/sha_core/n3718_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3620_187 )
);
defparam \top/processor/sha_core/n3620_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3620_s169  (
	.I0(\top/processor/sha_core/n3718_139 ),
	.I1(\top/processor/sha_core/n3718_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3620_189 )
);
defparam \top/processor/sha_core/n3620_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3620_s170  (
	.I0(\top/processor/sha_core/n3718_143 ),
	.I1(\top/processor/sha_core/n3718_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3620_191 )
);
defparam \top/processor/sha_core/n3620_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3620_s171  (
	.I0(\top/processor/sha_core/n3718_147 ),
	.I1(\top/processor/sha_core/n3718_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3620_193 )
);
defparam \top/processor/sha_core/n3620_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3621_s168  (
	.I0(\top/processor/sha_core/n3719_135 ),
	.I1(\top/processor/sha_core/n3719_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3621_187 )
);
defparam \top/processor/sha_core/n3621_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3621_s169  (
	.I0(\top/processor/sha_core/n3719_139 ),
	.I1(\top/processor/sha_core/n3719_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3621_189 )
);
defparam \top/processor/sha_core/n3621_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3621_s170  (
	.I0(\top/processor/sha_core/n3719_143 ),
	.I1(\top/processor/sha_core/n3719_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3621_191 )
);
defparam \top/processor/sha_core/n3621_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3621_s171  (
	.I0(\top/processor/sha_core/n3719_147 ),
	.I1(\top/processor/sha_core/n3719_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3621_193 )
);
defparam \top/processor/sha_core/n3621_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3622_s168  (
	.I0(\top/processor/sha_core/n3720_135 ),
	.I1(\top/processor/sha_core/n3720_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3622_187 )
);
defparam \top/processor/sha_core/n3622_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3622_s169  (
	.I0(\top/processor/sha_core/n3720_139 ),
	.I1(\top/processor/sha_core/n3720_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3622_189 )
);
defparam \top/processor/sha_core/n3622_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3622_s170  (
	.I0(\top/processor/sha_core/n3720_143 ),
	.I1(\top/processor/sha_core/n3720_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3622_191 )
);
defparam \top/processor/sha_core/n3622_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3622_s171  (
	.I0(\top/processor/sha_core/n3720_147 ),
	.I1(\top/processor/sha_core/n3720_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3622_193 )
);
defparam \top/processor/sha_core/n3622_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3623_s168  (
	.I0(\top/processor/sha_core/n3721_135 ),
	.I1(\top/processor/sha_core/n3721_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3623_187 )
);
defparam \top/processor/sha_core/n3623_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3623_s169  (
	.I0(\top/processor/sha_core/n3721_139 ),
	.I1(\top/processor/sha_core/n3721_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3623_189 )
);
defparam \top/processor/sha_core/n3623_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3623_s170  (
	.I0(\top/processor/sha_core/n3721_143 ),
	.I1(\top/processor/sha_core/n3721_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3623_191 )
);
defparam \top/processor/sha_core/n3623_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3623_s171  (
	.I0(\top/processor/sha_core/n3721_147 ),
	.I1(\top/processor/sha_core/n3721_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3623_193 )
);
defparam \top/processor/sha_core/n3623_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3624_s168  (
	.I0(\top/processor/sha_core/n3722_135 ),
	.I1(\top/processor/sha_core/n3722_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3624_187 )
);
defparam \top/processor/sha_core/n3624_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3624_s169  (
	.I0(\top/processor/sha_core/n3722_139 ),
	.I1(\top/processor/sha_core/n3722_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3624_189 )
);
defparam \top/processor/sha_core/n3624_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3624_s170  (
	.I0(\top/processor/sha_core/n3722_143 ),
	.I1(\top/processor/sha_core/n3722_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3624_191 )
);
defparam \top/processor/sha_core/n3624_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3624_s171  (
	.I0(\top/processor/sha_core/n3722_147 ),
	.I1(\top/processor/sha_core/n3722_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3624_193 )
);
defparam \top/processor/sha_core/n3624_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3625_s168  (
	.I0(\top/processor/sha_core/n3723_135 ),
	.I1(\top/processor/sha_core/n3723_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3625_187 )
);
defparam \top/processor/sha_core/n3625_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3625_s169  (
	.I0(\top/processor/sha_core/n3723_139 ),
	.I1(\top/processor/sha_core/n3723_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3625_189 )
);
defparam \top/processor/sha_core/n3625_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3625_s170  (
	.I0(\top/processor/sha_core/n3723_143 ),
	.I1(\top/processor/sha_core/n3723_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3625_191 )
);
defparam \top/processor/sha_core/n3625_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3625_s171  (
	.I0(\top/processor/sha_core/n3723_147 ),
	.I1(\top/processor/sha_core/n3723_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3625_193 )
);
defparam \top/processor/sha_core/n3625_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3626_s168  (
	.I0(\top/processor/sha_core/n3724_135 ),
	.I1(\top/processor/sha_core/n3724_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3626_187 )
);
defparam \top/processor/sha_core/n3626_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3626_s169  (
	.I0(\top/processor/sha_core/n3724_139 ),
	.I1(\top/processor/sha_core/n3724_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3626_189 )
);
defparam \top/processor/sha_core/n3626_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3626_s170  (
	.I0(\top/processor/sha_core/n3724_143 ),
	.I1(\top/processor/sha_core/n3724_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3626_191 )
);
defparam \top/processor/sha_core/n3626_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3626_s171  (
	.I0(\top/processor/sha_core/n3724_147 ),
	.I1(\top/processor/sha_core/n3724_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3626_193 )
);
defparam \top/processor/sha_core/n3626_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3627_s168  (
	.I0(\top/processor/sha_core/n3725_135 ),
	.I1(\top/processor/sha_core/n3725_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3627_187 )
);
defparam \top/processor/sha_core/n3627_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3627_s169  (
	.I0(\top/processor/sha_core/n3725_139 ),
	.I1(\top/processor/sha_core/n3725_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3627_189 )
);
defparam \top/processor/sha_core/n3627_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3627_s170  (
	.I0(\top/processor/sha_core/n3725_143 ),
	.I1(\top/processor/sha_core/n3725_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3627_191 )
);
defparam \top/processor/sha_core/n3627_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3627_s171  (
	.I0(\top/processor/sha_core/n3725_147 ),
	.I1(\top/processor/sha_core/n3725_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3627_193 )
);
defparam \top/processor/sha_core/n3627_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3628_s168  (
	.I0(\top/processor/sha_core/n3726_135 ),
	.I1(\top/processor/sha_core/n3726_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3628_187 )
);
defparam \top/processor/sha_core/n3628_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3628_s169  (
	.I0(\top/processor/sha_core/n3726_139 ),
	.I1(\top/processor/sha_core/n3726_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3628_189 )
);
defparam \top/processor/sha_core/n3628_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3628_s170  (
	.I0(\top/processor/sha_core/n3726_143 ),
	.I1(\top/processor/sha_core/n3726_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3628_191 )
);
defparam \top/processor/sha_core/n3628_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3628_s171  (
	.I0(\top/processor/sha_core/n3726_147 ),
	.I1(\top/processor/sha_core/n3726_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3628_193 )
);
defparam \top/processor/sha_core/n3628_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3629_s168  (
	.I0(\top/processor/sha_core/n3727_135 ),
	.I1(\top/processor/sha_core/n3727_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3629_187 )
);
defparam \top/processor/sha_core/n3629_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3629_s169  (
	.I0(\top/processor/sha_core/n3727_139 ),
	.I1(\top/processor/sha_core/n3727_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3629_189 )
);
defparam \top/processor/sha_core/n3629_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3629_s170  (
	.I0(\top/processor/sha_core/n3727_143 ),
	.I1(\top/processor/sha_core/n3727_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3629_191 )
);
defparam \top/processor/sha_core/n3629_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3629_s171  (
	.I0(\top/processor/sha_core/n3727_147 ),
	.I1(\top/processor/sha_core/n3727_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3629_193 )
);
defparam \top/processor/sha_core/n3629_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3630_s168  (
	.I0(\top/processor/sha_core/n3728_135 ),
	.I1(\top/processor/sha_core/n3728_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3630_187 )
);
defparam \top/processor/sha_core/n3630_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3630_s169  (
	.I0(\top/processor/sha_core/n3728_139 ),
	.I1(\top/processor/sha_core/n3728_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3630_189 )
);
defparam \top/processor/sha_core/n3630_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3630_s170  (
	.I0(\top/processor/sha_core/n3728_143 ),
	.I1(\top/processor/sha_core/n3728_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3630_191 )
);
defparam \top/processor/sha_core/n3630_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3630_s171  (
	.I0(\top/processor/sha_core/n3728_147 ),
	.I1(\top/processor/sha_core/n3728_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3630_193 )
);
defparam \top/processor/sha_core/n3630_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3631_s168  (
	.I0(\top/processor/sha_core/n3729_135 ),
	.I1(\top/processor/sha_core/n3729_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3631_187 )
);
defparam \top/processor/sha_core/n3631_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3631_s169  (
	.I0(\top/processor/sha_core/n3729_139 ),
	.I1(\top/processor/sha_core/n3729_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3631_189 )
);
defparam \top/processor/sha_core/n3631_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3631_s170  (
	.I0(\top/processor/sha_core/n3729_143 ),
	.I1(\top/processor/sha_core/n3729_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3631_191 )
);
defparam \top/processor/sha_core/n3631_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3631_s171  (
	.I0(\top/processor/sha_core/n3729_147 ),
	.I1(\top/processor/sha_core/n3729_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3631_193 )
);
defparam \top/processor/sha_core/n3631_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3632_s168  (
	.I0(\top/processor/sha_core/n3730_135 ),
	.I1(\top/processor/sha_core/n3730_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3632_187 )
);
defparam \top/processor/sha_core/n3632_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3632_s169  (
	.I0(\top/processor/sha_core/n3730_139 ),
	.I1(\top/processor/sha_core/n3730_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3632_189 )
);
defparam \top/processor/sha_core/n3632_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3632_s170  (
	.I0(\top/processor/sha_core/n3730_143 ),
	.I1(\top/processor/sha_core/n3730_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3632_191 )
);
defparam \top/processor/sha_core/n3632_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3632_s171  (
	.I0(\top/processor/sha_core/n3730_147 ),
	.I1(\top/processor/sha_core/n3730_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3632_193 )
);
defparam \top/processor/sha_core/n3632_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3633_s168  (
	.I0(\top/processor/sha_core/n3731_135 ),
	.I1(\top/processor/sha_core/n3731_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3633_187 )
);
defparam \top/processor/sha_core/n3633_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3633_s169  (
	.I0(\top/processor/sha_core/n3731_139 ),
	.I1(\top/processor/sha_core/n3731_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3633_189 )
);
defparam \top/processor/sha_core/n3633_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3633_s170  (
	.I0(\top/processor/sha_core/n3731_143 ),
	.I1(\top/processor/sha_core/n3731_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3633_191 )
);
defparam \top/processor/sha_core/n3633_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3633_s171  (
	.I0(\top/processor/sha_core/n3731_147 ),
	.I1(\top/processor/sha_core/n3731_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3633_193 )
);
defparam \top/processor/sha_core/n3633_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3634_s168  (
	.I0(\top/processor/sha_core/n3732_135 ),
	.I1(\top/processor/sha_core/n3732_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3634_187 )
);
defparam \top/processor/sha_core/n3634_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3634_s169  (
	.I0(\top/processor/sha_core/n3732_139 ),
	.I1(\top/processor/sha_core/n3732_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3634_189 )
);
defparam \top/processor/sha_core/n3634_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3634_s170  (
	.I0(\top/processor/sha_core/n3732_143 ),
	.I1(\top/processor/sha_core/n3732_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3634_191 )
);
defparam \top/processor/sha_core/n3634_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3634_s171  (
	.I0(\top/processor/sha_core/n3732_147 ),
	.I1(\top/processor/sha_core/n3732_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3634_193 )
);
defparam \top/processor/sha_core/n3634_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3635_s168  (
	.I0(\top/processor/sha_core/n3733_135 ),
	.I1(\top/processor/sha_core/n3733_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3635_187 )
);
defparam \top/processor/sha_core/n3635_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3635_s169  (
	.I0(\top/processor/sha_core/n3733_139 ),
	.I1(\top/processor/sha_core/n3733_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3635_189 )
);
defparam \top/processor/sha_core/n3635_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3635_s170  (
	.I0(\top/processor/sha_core/n3733_143 ),
	.I1(\top/processor/sha_core/n3733_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3635_191 )
);
defparam \top/processor/sha_core/n3635_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3635_s171  (
	.I0(\top/processor/sha_core/n3733_147 ),
	.I1(\top/processor/sha_core/n3733_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3635_193 )
);
defparam \top/processor/sha_core/n3635_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3636_s168  (
	.I0(\top/processor/sha_core/n3734_135 ),
	.I1(\top/processor/sha_core/n3734_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3636_187 )
);
defparam \top/processor/sha_core/n3636_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3636_s169  (
	.I0(\top/processor/sha_core/n3734_139 ),
	.I1(\top/processor/sha_core/n3734_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3636_189 )
);
defparam \top/processor/sha_core/n3636_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3636_s170  (
	.I0(\top/processor/sha_core/n3734_143 ),
	.I1(\top/processor/sha_core/n3734_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3636_191 )
);
defparam \top/processor/sha_core/n3636_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3636_s171  (
	.I0(\top/processor/sha_core/n3734_147 ),
	.I1(\top/processor/sha_core/n3734_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3636_193 )
);
defparam \top/processor/sha_core/n3636_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3637_s168  (
	.I0(\top/processor/sha_core/n3735_135 ),
	.I1(\top/processor/sha_core/n3735_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3637_187 )
);
defparam \top/processor/sha_core/n3637_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3637_s169  (
	.I0(\top/processor/sha_core/n3735_139 ),
	.I1(\top/processor/sha_core/n3735_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3637_189 )
);
defparam \top/processor/sha_core/n3637_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3637_s170  (
	.I0(\top/processor/sha_core/n3735_143 ),
	.I1(\top/processor/sha_core/n3735_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3637_191 )
);
defparam \top/processor/sha_core/n3637_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3637_s171  (
	.I0(\top/processor/sha_core/n3735_147 ),
	.I1(\top/processor/sha_core/n3735_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3637_193 )
);
defparam \top/processor/sha_core/n3637_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3638_s168  (
	.I0(\top/processor/sha_core/n3736_135 ),
	.I1(\top/processor/sha_core/n3736_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3638_187 )
);
defparam \top/processor/sha_core/n3638_s168 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3638_s169  (
	.I0(\top/processor/sha_core/n3736_139 ),
	.I1(\top/processor/sha_core/n3736_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3638_189 )
);
defparam \top/processor/sha_core/n3638_s169 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3638_s170  (
	.I0(\top/processor/sha_core/n3736_143 ),
	.I1(\top/processor/sha_core/n3736_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3638_191 )
);
defparam \top/processor/sha_core/n3638_s170 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3638_s171  (
	.I0(\top/processor/sha_core/n3736_147 ),
	.I1(\top/processor/sha_core/n3736_145 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n3638_193 )
);
defparam \top/processor/sha_core/n3638_s171 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n293_s5621  (
	.I0(\top/processor/sha_core/n293_7225 ),
	.I1(\top/processor/sha_core/n293_7226 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7162 )
);
defparam \top/processor/sha_core/n293_s5621 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n293_s5622  (
	.I0(\top/processor/sha_core/n293_7227 ),
	.I1(\top/processor/sha_core/n293_7228 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7164 )
);
defparam \top/processor/sha_core/n293_s5622 .INIT=8'h35;
LUT4 \top/processor/sha_core/n293_s5623  (
	.I0(\top/processor/sha_core/n293_7229 ),
	.I1(\top/processor/sha_core/n293_7230 ),
	.I2(\top/processor/sha_core/n293_7231 ),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7166 )
);
defparam \top/processor/sha_core/n293_s5623 .INIT=16'h0B0C;
LUT3 \top/processor/sha_core/n293_s5624  (
	.I0(\top/processor/sha_core/n293_7232 ),
	.I1(\top/processor/sha_core/n293_7233 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7168 )
);
defparam \top/processor/sha_core/n293_s5624 .INIT=8'h35;
LUT4 \top/processor/sha_core/n293_s5625  (
	.I0(\top/processor/sha_core/n293_7386 ),
	.I1(\top/processor/sha_core/n293_7235 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7236 ),
	.F(\top/processor/sha_core/n293_7170 )
);
defparam \top/processor/sha_core/n293_s5625 .INIT=16'hCFA0;
LUT3 \top/processor/sha_core/n293_s5626  (
	.I0(\top/processor/sha_core/n293_7237 ),
	.I1(\top/processor/sha_core/n293_7238 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7172 )
);
defparam \top/processor/sha_core/n293_s5626 .INIT=8'h3A;
LUT3 \top/processor/sha_core/n293_s5627  (
	.I0(\top/processor/sha_core/n293_7239 ),
	.I1(\top/processor/sha_core/n293_7240 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7174 )
);
defparam \top/processor/sha_core/n293_s5627 .INIT=8'hCA;
LUT4 \top/processor/sha_core/n293_s5628  (
	.I0(\top/processor/sha_core/n293_7241 ),
	.I1(\top/processor/sha_core/n293_7242 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7243 ),
	.F(\top/processor/sha_core/n293_7176 )
);
defparam \top/processor/sha_core/n293_s5628 .INIT=16'hA03F;
LUT4 \top/processor/sha_core/n293_s5629  (
	.I0(\top/processor/sha_core/n293_7244 ),
	.I1(\top/processor/sha_core/n293_7245 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7246 ),
	.F(\top/processor/sha_core/n293_7178 )
);
defparam \top/processor/sha_core/n293_s5629 .INIT=16'h3FA0;
LUT3 \top/processor/sha_core/n293_s5630  (
	.I0(\top/processor/sha_core/n293_7247 ),
	.I1(\top/processor/sha_core/n293_7248 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7180 )
);
defparam \top/processor/sha_core/n293_s5630 .INIT=8'h3A;
LUT4 \top/processor/sha_core/n293_s5631  (
	.I0(\top/processor/sha_core/n293_7249 ),
	.I1(\top/processor/sha_core/n293_7250 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7251 ),
	.F(\top/processor/sha_core/n293_7182 )
);
defparam \top/processor/sha_core/n293_s5631 .INIT=16'h3F50;
LUT4 \top/processor/sha_core/n293_s5632  (
	.I0(\top/processor/sha_core/t [0]),
	.I1(\top/processor/sha_core/n293_7252 ),
	.I2(\top/processor/sha_core/n293_7253 ),
	.I3(\top/processor/sha_core/n293_7254 ),
	.F(\top/processor/sha_core/n293_7184 )
);
defparam \top/processor/sha_core/n293_s5632 .INIT=16'h7A70;
LUT4 \top/processor/sha_core/n293_s5633  (
	.I0(\top/processor/sha_core/n293_7255 ),
	.I1(\top/processor/sha_core/n293_7256 ),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/n293_7257 ),
	.F(\top/processor/sha_core/n293_7186 )
);
defparam \top/processor/sha_core/n293_s5633 .INIT=16'h3F50;
LUT4 \top/processor/sha_core/n293_s5634  (
	.I0(\top/processor/sha_core/n293_7258 ),
	.I1(\top/processor/sha_core/n293_7259 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7260 ),
	.F(\top/processor/sha_core/n293_7188 )
);
defparam \top/processor/sha_core/n293_s5634 .INIT=16'h503F;
LUT4 \top/processor/sha_core/n293_s5635  (
	.I0(\top/processor/sha_core/n293_7261 ),
	.I1(\top/processor/sha_core/n293_7262 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7263 ),
	.F(\top/processor/sha_core/n293_7190 )
);
defparam \top/processor/sha_core/n293_s5635 .INIT=16'h503F;
LUT4 \top/processor/sha_core/n293_s5636  (
	.I0(\top/processor/sha_core/n293_7264 ),
	.I1(\top/processor/sha_core/n293_7265 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7266 ),
	.F(\top/processor/sha_core/n293_7192 )
);
defparam \top/processor/sha_core/n293_s5636 .INIT=16'h3F50;
LUT3 \top/processor/sha_core/n293_s5637  (
	.I0(\top/processor/sha_core/n293_7267 ),
	.I1(\top/processor/sha_core/n293_7268 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7194 )
);
defparam \top/processor/sha_core/n293_s5637 .INIT=8'hCA;
LUT3 \top/processor/sha_core/n293_s5638  (
	.I0(\top/processor/sha_core/n293_7269 ),
	.I1(\top/processor/sha_core/n293_7270 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7196 )
);
defparam \top/processor/sha_core/n293_s5638 .INIT=8'hC5;
LUT4 \top/processor/sha_core/n293_s5639  (
	.I0(\top/processor/sha_core/n293_7271 ),
	.I1(\top/processor/sha_core/n293_7272 ),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/n293_7273 ),
	.F(\top/processor/sha_core/n293_7198 )
);
defparam \top/processor/sha_core/n293_s5639 .INIT=16'h3B38;
LUT4 \top/processor/sha_core/n293_s5640  (
	.I0(\top/processor/sha_core/n293_7274 ),
	.I1(\top/processor/sha_core/n293_7275 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7276 ),
	.F(\top/processor/sha_core/n293_7200 )
);
defparam \top/processor/sha_core/n293_s5640 .INIT=16'h50CF;
LUT4 \top/processor/sha_core/n293_s5641  (
	.I0(\top/processor/sha_core/n293_7277 ),
	.I1(\top/processor/sha_core/n293_7278 ),
	.I2(\top/processor/sha_core/n293_7279 ),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7202 )
);
defparam \top/processor/sha_core/n293_s5641 .INIT=16'h33E0;
LUT4 \top/processor/sha_core/n293_s5642  (
	.I0(\top/processor/sha_core/n293_7280 ),
	.I1(\top/processor/sha_core/n293_7281 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7282 ),
	.F(\top/processor/sha_core/n293_7204 )
);
defparam \top/processor/sha_core/n293_s5642 .INIT=16'hCF50;
LUT4 \top/processor/sha_core/n293_s5643  (
	.I0(\top/processor/sha_core/n293_7283 ),
	.I1(\top/processor/sha_core/n293_7284 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7285 ),
	.F(\top/processor/sha_core/n293_7206 )
);
defparam \top/processor/sha_core/n293_s5643 .INIT=16'hA0CF;
LUT3 \top/processor/sha_core/n293_s5644  (
	.I0(\top/processor/sha_core/n293_7286 ),
	.I1(\top/processor/sha_core/n293_7287 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7208 )
);
defparam \top/processor/sha_core/n293_s5644 .INIT=8'hC5;
LUT3 \top/processor/sha_core/n293_s5645  (
	.I0(\top/processor/sha_core/n293_7288 ),
	.I1(\top/processor/sha_core/n293_7289 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7210 )
);
defparam \top/processor/sha_core/n293_s5645 .INIT=8'hCA;
LUT4 \top/processor/sha_core/n293_s5646  (
	.I0(\top/processor/sha_core/n293_7290 ),
	.I1(\top/processor/sha_core/n293_7291 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7292 ),
	.F(\top/processor/sha_core/n293_7212 )
);
defparam \top/processor/sha_core/n293_s5646 .INIT=16'h3F50;
LUT4 \top/processor/sha_core/n293_s5647  (
	.I0(\top/processor/sha_core/n293_7293 ),
	.I1(\top/processor/sha_core/n293_7294 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7295 ),
	.F(\top/processor/sha_core/n293_7214 )
);
defparam \top/processor/sha_core/n293_s5647 .INIT=16'hCFA0;
LUT4 \top/processor/sha_core/n293_s5648  (
	.I0(\top/processor/sha_core/n293_7296 ),
	.I1(\top/processor/sha_core/n293_7297 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7298 ),
	.F(\top/processor/sha_core/n293_7216 )
);
defparam \top/processor/sha_core/n293_s5648 .INIT=16'hCF50;
LUT3 \top/processor/sha_core/n293_s5649  (
	.I0(\top/processor/sha_core/n293_7299 ),
	.I1(\top/processor/sha_core/n293_7300 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7218 )
);
defparam \top/processor/sha_core/n293_s5649 .INIT=8'h35;
LUT3 \top/processor/sha_core/n293_s5650  (
	.I0(\top/processor/sha_core/n293_7301 ),
	.I1(\top/processor/sha_core/n293_7302 ),
	.I2(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7220 )
);
defparam \top/processor/sha_core/n293_s5650 .INIT=8'h35;
LUT4 \top/processor/sha_core/n293_s5651  (
	.I0(\top/processor/sha_core/n293_7303 ),
	.I1(\top/processor/sha_core/n293_7304 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7305 ),
	.F(\top/processor/sha_core/n293_7222 )
);
defparam \top/processor/sha_core/n293_s5651 .INIT=16'h3D31;
LUT4 \top/processor/sha_core/n293_s5652  (
	.I0(\top/processor/sha_core/n293_7306 ),
	.I1(\top/processor/sha_core/n293_7307 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/n293_7308 ),
	.F(\top/processor/sha_core/n293_7224 )
);
defparam \top/processor/sha_core/n293_s5652 .INIT=16'hCF50;
LUT2 \top/processor/sha_core/n14445_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/n14445_10 )
);
defparam \top/processor/sha_core/n14445_s5 .INIT=4'h4;
LUT2 \top/processor/sha_core/n14442_s4  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/n3607_196 ),
	.F(\top/processor/sha_core/n14442_9 )
);
defparam \top/processor/sha_core/n14442_s4 .INIT=4'h2;
LUT4 \top/processor/sha_core/n14440_s4  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/w[31]_31_11 ),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.I3(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/n14440_9 )
);
defparam \top/processor/sha_core/n14440_s4 .INIT=16'h7800;
LUT3 \top/processor/sha_core/n14439_s4  (
	.I0(\top/processor/sha_core/n14439_10 ),
	.I1(\top/processor/sha_core/msg_idx [6]),
	.I2(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/n14439_9 )
);
defparam \top/processor/sha_core/n14439_s4 .INIT=8'h60;
LUT2 \top/processor/sha_core/n12134_s6  (
	.I0(\top/processor/sha_core/t [0]),
	.I1(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12134_11 )
);
defparam \top/processor/sha_core/n12134_s6 .INIT=4'h4;
LUT3 \top/processor/sha_core/n12133_s6  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [0]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12133_11 )
);
defparam \top/processor/sha_core/n12133_s6 .INIT=8'h60;
LUT4 \top/processor/sha_core/n12132_s6  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [0]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12132_11 )
);
defparam \top/processor/sha_core/n12132_s6 .INIT=16'h7800;
LUT3 \top/processor/sha_core/n12131_s6  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/n12131_12 ),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12131_11 )
);
defparam \top/processor/sha_core/n12131_s6 .INIT=8'h60;
LUT4 \top/processor/sha_core/n12130_s6  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/n12131_12 ),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12130_11 )
);
defparam \top/processor/sha_core/n12130_s6 .INIT=16'h7800;
LUT3 \top/processor/sha_core/n12129_s6  (
	.I0(\top/processor/sha_core/n12129_12 ),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12129_11 )
);
defparam \top/processor/sha_core/n12129_s6 .INIT=8'h60;
LUT3 \top/processor/sha_core/n12128_s6  (
	.I0(\top/processor/sha_core/n12128_12 ),
	.I1(\top/processor/sha_core/t [6]),
	.I2(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n12128_11 )
);
defparam \top/processor/sha_core/n12128_s6 .INIT=8'h60;
LUT2 \top/processor/sha_core/n3462_s4  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.F(\top/processor/sha_core/n3462_11 )
);
defparam \top/processor/sha_core/n3462_s4 .INIT=4'h9;
LUT3 \top/processor/sha_core/n3461_s4  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.F(\top/processor/sha_core/n3461_11 )
);
defparam \top/processor/sha_core/n3461_s4 .INIT=8'hE1;
LUT4 \top/processor/sha_core/n3460_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/msg_idx [4]),
	.F(\top/processor/sha_core/n3460_11 )
);
defparam \top/processor/sha_core/n3460_s4 .INIT=16'hFE01;
LUT4 \top/processor/sha_core/n3459_s3  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/w[0]_31_9 ),
	.I3(\top/processor/sha_core/msg_idx [5]),
	.F(\top/processor/sha_core/n3459_9 )
);
defparam \top/processor/sha_core/n3459_s3 .INIT=16'hEF10;
LUT3 \top/processor/sha_core/n3578_s4  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/n3578_12 ),
	.I2(\top/processor/sha_core/msg_idx [4]),
	.F(\top/processor/sha_core/n3578_11 )
);
defparam \top/processor/sha_core/n3578_s4 .INIT=8'hE1;
LUT2 \top/processor/sha_core/n3834_s3  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.F(\top/processor/sha_core/n3834_9 )
);
defparam \top/processor/sha_core/n3834_s3 .INIT=4'h9;
LUT3 \top/processor/sha_core/n3766_s1  (
	.I0(\top/processor/sha_core/n3766_6 ),
	.I1(\top/processor/sha_core/n3766_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3766_4 )
);
defparam \top/processor/sha_core/n3766_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3766_s2  (
	.I0(\top/processor/sha_core/n3766_9 ),
	.I1(\top/processor/sha_core/n3766_10 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3766_5 )
);
defparam \top/processor/sha_core/n3766_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3767_s1  (
	.I0(\top/processor/sha_core/n3767_6 ),
	.I1(\top/processor/sha_core/n3767_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3767_4 )
);
defparam \top/processor/sha_core/n3767_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3767_s2  (
	.I0(\top/processor/sha_core/n3767_8 ),
	.I1(\top/processor/sha_core/n3767_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3767_5 )
);
defparam \top/processor/sha_core/n3767_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3768_s1  (
	.I0(\top/processor/sha_core/n3768_6 ),
	.I1(\top/processor/sha_core/n3768_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3768_4 )
);
defparam \top/processor/sha_core/n3768_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3768_s2  (
	.I0(\top/processor/sha_core/n3768_8 ),
	.I1(\top/processor/sha_core/n3768_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3768_5 )
);
defparam \top/processor/sha_core/n3768_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3769_s1  (
	.I0(\top/processor/sha_core/n3769_7 ),
	.I1(\top/processor/sha_core/n3769_8 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3769_4 )
);
defparam \top/processor/sha_core/n3769_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3769_s2  (
	.I0(\top/processor/sha_core/n3769_9 ),
	.I1(\top/processor/sha_core/n3769_10 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3769_5 )
);
defparam \top/processor/sha_core/n3769_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3769_s3  (
	.I0(\top/processor/sha_core/n3769_11 ),
	.I1(\top/processor/sha_core/n3769_12 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3769_6 )
);
defparam \top/processor/sha_core/n3769_s3 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3770_s1  (
	.I0(\top/processor/sha_core/n3770_6 ),
	.I1(\top/processor/sha_core/n3770_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3770_4 )
);
defparam \top/processor/sha_core/n3770_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3770_s2  (
	.I0(\top/processor/sha_core/n3770_8 ),
	.I1(\top/processor/sha_core/n3770_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3770_5 )
);
defparam \top/processor/sha_core/n3770_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3771_s1  (
	.I0(\top/processor/sha_core/n3771_6 ),
	.I1(\top/processor/sha_core/n3771_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3771_4 )
);
defparam \top/processor/sha_core/n3771_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3771_s2  (
	.I0(\top/processor/sha_core/n3771_8 ),
	.I1(\top/processor/sha_core/n3771_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3771_5 )
);
defparam \top/processor/sha_core/n3771_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3772_s1  (
	.I0(\top/processor/sha_core/n3772_6 ),
	.I1(\top/processor/sha_core/n3772_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3772_4 )
);
defparam \top/processor/sha_core/n3772_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3772_s2  (
	.I0(\top/processor/sha_core/n3772_8 ),
	.I1(\top/processor/sha_core/n3772_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3772_5 )
);
defparam \top/processor/sha_core/n3772_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3773_s1  (
	.I0(\top/processor/sha_core/n3773_6 ),
	.I1(\top/processor/sha_core/n3773_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3773_4 )
);
defparam \top/processor/sha_core/n3773_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3773_s2  (
	.I0(\top/processor/sha_core/n3773_8 ),
	.I1(\top/processor/sha_core/n3773_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3773_5 )
);
defparam \top/processor/sha_core/n3773_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3774_s1  (
	.I0(\top/processor/sha_core/n3774_6 ),
	.I1(\top/processor/sha_core/n3774_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3774_4 )
);
defparam \top/processor/sha_core/n3774_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3774_s2  (
	.I0(\top/processor/sha_core/n3774_8 ),
	.I1(\top/processor/sha_core/n3774_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3774_5 )
);
defparam \top/processor/sha_core/n3774_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3775_s1  (
	.I0(\top/processor/sha_core/n3775_6 ),
	.I1(\top/processor/sha_core/n3775_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3775_4 )
);
defparam \top/processor/sha_core/n3775_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3775_s2  (
	.I0(\top/processor/sha_core/n3775_8 ),
	.I1(\top/processor/sha_core/n3775_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3775_5 )
);
defparam \top/processor/sha_core/n3775_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3776_s1  (
	.I0(\top/processor/sha_core/n3776_6 ),
	.I1(\top/processor/sha_core/n3776_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3776_4 )
);
defparam \top/processor/sha_core/n3776_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3776_s2  (
	.I0(\top/processor/sha_core/n3776_8 ),
	.I1(\top/processor/sha_core/n3776_9 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3776_5 )
);
defparam \top/processor/sha_core/n3776_s2 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3777_s1  (
	.I0(\top/processor/sha_core/n3777_5 ),
	.I1(\top/processor/sha_core/n3777_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3777_4 )
);
defparam \top/processor/sha_core/n3777_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3778_s1  (
	.I0(\top/processor/sha_core/n3778_5 ),
	.I1(\top/processor/sha_core/n3778_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3778_4 )
);
defparam \top/processor/sha_core/n3778_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3779_s1  (
	.I0(\top/processor/sha_core/n3779_5 ),
	.I1(\top/processor/sha_core/n3779_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3779_4 )
);
defparam \top/processor/sha_core/n3779_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3780_s1  (
	.I0(\top/processor/sha_core/n3780_5 ),
	.I1(\top/processor/sha_core/n3780_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3780_4 )
);
defparam \top/processor/sha_core/n3780_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3781_s1  (
	.I0(\top/processor/sha_core/n3781_5 ),
	.I1(\top/processor/sha_core/n3781_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3781_4 )
);
defparam \top/processor/sha_core/n3781_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3782_s1  (
	.I0(\top/processor/sha_core/n3782_5 ),
	.I1(\top/processor/sha_core/n3782_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3782_4 )
);
defparam \top/processor/sha_core/n3782_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3783_s1  (
	.I0(\top/processor/sha_core/n3783_5 ),
	.I1(\top/processor/sha_core/n3783_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3783_4 )
);
defparam \top/processor/sha_core/n3783_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3784_s1  (
	.I0(\top/processor/sha_core/n3784_5 ),
	.I1(\top/processor/sha_core/n3784_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3784_4 )
);
defparam \top/processor/sha_core/n3784_s1 .INIT=8'hAC;
LUT3 \top/processor/sha_core/n3785_s1  (
	.I0(\top/processor/sha_core/n3785_5 ),
	.I1(\top/processor/sha_core/n3785_6 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.F(\top/processor/sha_core/n3785_4 )
);
defparam \top/processor/sha_core/n3785_s1 .INIT=8'hAC;
LUT4 \top/processor/sha_core/n8430_s1  (
	.I0(\top/processor/sha_core/n8430_7 ),
	.I1(\top/processor/sha_core/n8430_8 ),
	.I2(\top/processor/sha_core/n8430_9 ),
	.I3(\top/processor/sha_core/n8430_10 ),
	.F(\top/processor/sha_core/n8430_4 )
);
defparam \top/processor/sha_core/n8430_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8430_s2  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [511]),
	.I2(\top/processor/sha_core/n8430_12 ),
	.I3(\top/processor/sha_core/n8430_13 ),
	.F(\top/processor/sha_core/n8430_5 )
);
defparam \top/processor/sha_core/n8430_s2 .INIT=16'h7000;
LUT3 \top/processor/sha_core/n8430_s3  (
	.I0(\top/processor/sha_core/msg_idx [6]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.F(\top/processor/sha_core/n8430_6 )
);
defparam \top/processor/sha_core/n8430_s3 .INIT=8'h01;
LUT4 \top/processor/sha_core/n8431_s1  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [478]),
	.I2(\top/processor/sha_core/n8431_7 ),
	.I3(\top/processor/sha_core/n8431_8 ),
	.F(\top/processor/sha_core/n8431_4 )
);
defparam \top/processor/sha_core/n8431_s1 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8431_s2  (
	.I0(\top/processor/sha_core/n8431_9 ),
	.I1(\top/processor/sha_core/n8431_10 ),
	.I2(\top/processor/sha_core/n8431_11 ),
	.I3(\top/processor/sha_core/n8431_12 ),
	.F(\top/processor/sha_core/n8431_5 )
);
defparam \top/processor/sha_core/n8431_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8432_s1  (
	.I0(\top/processor/sha_core/n8432_6 ),
	.I1(\top/processor/sha_core/n8432_7 ),
	.I2(\top/processor/sha_core/n8432_8 ),
	.I3(\top/processor/sha_core/n8432_9 ),
	.F(\top/processor/sha_core/n8432_4 )
);
defparam \top/processor/sha_core/n8432_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8432_s2  (
	.I0(\top/processor/sha_core/w[3]_31_9 ),
	.I1(\top/processor/core_block [413]),
	.I2(\top/processor/sha_core/n8432_10 ),
	.I3(\top/processor/sha_core/n8432_11 ),
	.F(\top/processor/sha_core/n8432_5 )
);
defparam \top/processor/sha_core/n8432_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8433_s1  (
	.I0(\top/processor/sha_core/n8433_6 ),
	.I1(\top/processor/sha_core/n8433_7 ),
	.I2(\top/processor/sha_core/n8433_8 ),
	.I3(\top/processor/sha_core/n8433_9 ),
	.F(\top/processor/sha_core/n8433_4 )
);
defparam \top/processor/sha_core/n8433_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8433_s2  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [188]),
	.I2(\top/processor/sha_core/n8433_10 ),
	.I3(\top/processor/sha_core/n8433_11 ),
	.F(\top/processor/sha_core/n8433_5 )
);
defparam \top/processor/sha_core/n8433_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8434_s1  (
	.I0(\top/processor/sha_core/n8434_6 ),
	.I1(\top/processor/sha_core/n8434_7 ),
	.I2(\top/processor/sha_core/n8434_8 ),
	.I3(\top/processor/sha_core/n8434_9 ),
	.F(\top/processor/sha_core/n8434_4 )
);
defparam \top/processor/sha_core/n8434_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8434_s2  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [187]),
	.I2(\top/processor/sha_core/n8434_10 ),
	.I3(\top/processor/sha_core/n8434_11 ),
	.F(\top/processor/sha_core/n8434_5 )
);
defparam \top/processor/sha_core/n8434_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8435_s1  (
	.I0(\top/processor/sha_core/n8435_6 ),
	.I1(\top/processor/sha_core/n8435_7 ),
	.I2(\top/processor/sha_core/n8435_8 ),
	.I3(\top/processor/sha_core/n8435_9 ),
	.F(\top/processor/sha_core/n8435_4 )
);
defparam \top/processor/sha_core/n8435_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8435_s2  (
	.I0(\top/processor/sha_core/n8435_10 ),
	.I1(\top/processor/sha_core/n8435_11 ),
	.I2(\top/processor/sha_core/n8435_12 ),
	.I3(\top/processor/sha_core/n8435_13 ),
	.F(\top/processor/sha_core/n8435_5 )
);
defparam \top/processor/sha_core/n8435_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8436_s1  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [121]),
	.I2(\top/processor/sha_core/n8436_6 ),
	.I3(\top/processor/sha_core/n8436_7 ),
	.F(\top/processor/sha_core/n8436_4 )
);
defparam \top/processor/sha_core/n8436_s1 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8436_s2  (
	.I0(\top/processor/sha_core/n8436_8 ),
	.I1(\top/processor/sha_core/n8436_9 ),
	.I2(\top/processor/sha_core/n8436_10 ),
	.I3(\top/processor/sha_core/n8436_11 ),
	.F(\top/processor/sha_core/n8436_5 )
);
defparam \top/processor/sha_core/n8436_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8437_s1  (
	.I0(\top/processor/sha_core/n8437_6 ),
	.I1(\top/processor/sha_core/n8437_7 ),
	.I2(\top/processor/sha_core/n8437_8 ),
	.I3(\top/processor/sha_core/n8437_9 ),
	.F(\top/processor/sha_core/n8437_4 )
);
defparam \top/processor/sha_core/n8437_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8437_s2  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [184]),
	.I2(\top/processor/sha_core/n8437_10 ),
	.I3(\top/processor/sha_core/n8437_11 ),
	.F(\top/processor/sha_core/n8437_5 )
);
defparam \top/processor/sha_core/n8437_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8438_s1  (
	.I0(\top/processor/sha_core/n8438_6 ),
	.I1(\top/processor/sha_core/n8438_7 ),
	.I2(\top/processor/sha_core/n8438_8 ),
	.I3(\top/processor/sha_core/n8438_9 ),
	.F(\top/processor/sha_core/n8438_4 )
);
defparam \top/processor/sha_core/n8438_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8438_s2  (
	.I0(\top/processor/sha_core/w[14]_31_9 ),
	.I1(\top/processor/core_block [55]),
	.I2(\top/processor/sha_core/n8438_10 ),
	.I3(\top/processor/sha_core/n8438_11 ),
	.F(\top/processor/sha_core/n8438_5 )
);
defparam \top/processor/sha_core/n8438_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8439_s1  (
	.I0(\top/processor/sha_core/w[3]_31_9 ),
	.I1(\top/processor/core_block [406]),
	.I2(\top/processor/sha_core/n8439_5 ),
	.I3(\top/processor/sha_core/n8439_6 ),
	.F(\top/processor/sha_core/n8439_4 )
);
defparam \top/processor/sha_core/n8439_s1 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8440_s1  (
	.I0(\top/processor/sha_core/n8440_6 ),
	.I1(\top/processor/sha_core/n8440_7 ),
	.I2(\top/processor/sha_core/n8440_8 ),
	.I3(\top/processor/sha_core/n8440_9 ),
	.F(\top/processor/sha_core/n8440_4 )
);
defparam \top/processor/sha_core/n8440_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8440_s2  (
	.I0(\top/processor/sha_core/w[3]_31_9 ),
	.I1(\top/processor/core_block [405]),
	.I2(\top/processor/sha_core/n8440_10 ),
	.I3(\top/processor/sha_core/n8440_11 ),
	.F(\top/processor/sha_core/n8440_5 )
);
defparam \top/processor/sha_core/n8440_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8441_s1  (
	.I0(\top/processor/sha_core/n8441_6 ),
	.I1(\top/processor/sha_core/n8441_7 ),
	.I2(\top/processor/sha_core/n8441_8 ),
	.I3(\top/processor/sha_core/n8441_9 ),
	.F(\top/processor/sha_core/n8441_4 )
);
defparam \top/processor/sha_core/n8441_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8441_s2  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [500]),
	.I2(\top/processor/sha_core/n8441_10 ),
	.I3(\top/processor/sha_core/n8441_11 ),
	.F(\top/processor/sha_core/n8441_5 )
);
defparam \top/processor/sha_core/n8441_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8442_s1  (
	.I0(\top/processor/sha_core/n8442_5 ),
	.I1(\top/processor/sha_core/n8442_6 ),
	.I2(\top/processor/sha_core/n8442_7 ),
	.I3(\top/processor/sha_core/n8442_8 ),
	.F(\top/processor/sha_core/n8442_4 )
);
defparam \top/processor/sha_core/n8442_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8443_s1  (
	.I0(\top/processor/sha_core/n8443_6 ),
	.I1(\top/processor/sha_core/n8443_7 ),
	.I2(\top/processor/sha_core/n8443_8 ),
	.I3(\top/processor/sha_core/n8443_9 ),
	.F(\top/processor/sha_core/n8443_4 )
);
defparam \top/processor/sha_core/n8443_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8443_s2  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [306]),
	.I2(\top/processor/sha_core/n8443_10 ),
	.I3(\top/processor/sha_core/n8443_11 ),
	.F(\top/processor/sha_core/n8443_5 )
);
defparam \top/processor/sha_core/n8443_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8444_s1  (
	.I0(\top/processor/sha_core/n8444_6 ),
	.I1(\top/processor/sha_core/n8444_7 ),
	.I2(\top/processor/sha_core/n8444_8 ),
	.I3(\top/processor/sha_core/n8444_9 ),
	.F(\top/processor/sha_core/n8444_4 )
);
defparam \top/processor/sha_core/n8444_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8444_s2  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/core_block [241]),
	.I2(\top/processor/sha_core/n8444_10 ),
	.I3(\top/processor/sha_core/n8444_11 ),
	.F(\top/processor/sha_core/n8444_5 )
);
defparam \top/processor/sha_core/n8444_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8445_s1  (
	.I0(\top/processor/sha_core/n8445_6 ),
	.I1(\top/processor/sha_core/n8445_7 ),
	.I2(\top/processor/sha_core/n8445_8 ),
	.I3(\top/processor/sha_core/n8445_9 ),
	.F(\top/processor/sha_core/n8445_4 )
);
defparam \top/processor/sha_core/n8445_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8445_s2  (
	.I0(\top/processor/sha_core/n8445_10 ),
	.I1(\top/processor/sha_core/n8445_11 ),
	.I2(\top/processor/sha_core/n8445_12 ),
	.I3(\top/processor/sha_core/n8445_13 ),
	.F(\top/processor/sha_core/n8445_5 )
);
defparam \top/processor/sha_core/n8445_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8446_s1  (
	.I0(\top/processor/sha_core/n8446_6 ),
	.I1(\top/processor/sha_core/n8446_7 ),
	.I2(\top/processor/sha_core/n8446_8 ),
	.I3(\top/processor/sha_core/n8446_9 ),
	.F(\top/processor/sha_core/n8446_4 )
);
defparam \top/processor/sha_core/n8446_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8446_s2  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [175]),
	.I2(\top/processor/sha_core/n8446_10 ),
	.I3(\top/processor/sha_core/n8446_11 ),
	.F(\top/processor/sha_core/n8446_5 )
);
defparam \top/processor/sha_core/n8446_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8447_s1  (
	.I0(\top/processor/sha_core/n8447_6 ),
	.I1(\top/processor/sha_core/n8447_7 ),
	.I2(\top/processor/sha_core/n8447_8 ),
	.I3(\top/processor/sha_core/n8447_9 ),
	.F(\top/processor/sha_core/n8447_4 )
);
defparam \top/processor/sha_core/n8447_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8447_s2  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [206]),
	.I2(\top/processor/sha_core/n8447_10 ),
	.I3(\top/processor/sha_core/n8447_11 ),
	.F(\top/processor/sha_core/n8447_5 )
);
defparam \top/processor/sha_core/n8447_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8448_s1  (
	.I0(\top/processor/sha_core/n8448_6 ),
	.I1(\top/processor/sha_core/n8448_7 ),
	.I2(\top/processor/sha_core/n8448_8 ),
	.I3(\top/processor/sha_core/n8448_9 ),
	.F(\top/processor/sha_core/n8448_4 )
);
defparam \top/processor/sha_core/n8448_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8448_s2  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [493]),
	.I2(\top/processor/sha_core/n8448_10 ),
	.I3(\top/processor/sha_core/n8448_11 ),
	.F(\top/processor/sha_core/n8448_5 )
);
defparam \top/processor/sha_core/n8448_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8449_s1  (
	.I0(\top/processor/sha_core/n8449_6 ),
	.I1(\top/processor/sha_core/n8449_7 ),
	.I2(\top/processor/sha_core/n8449_8 ),
	.I3(\top/processor/sha_core/n8449_9 ),
	.F(\top/processor/sha_core/n8449_4 )
);
defparam \top/processor/sha_core/n8449_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8449_s2  (
	.I0(\top/processor/sha_core/w[14]_31_9 ),
	.I1(\top/processor/core_block [44]),
	.I2(\top/processor/sha_core/n8449_10 ),
	.I3(\top/processor/sha_core/n8449_11 ),
	.F(\top/processor/sha_core/n8449_5 )
);
defparam \top/processor/sha_core/n8449_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8450_s1  (
	.I0(\top/processor/sha_core/n8450_5 ),
	.I1(\top/processor/sha_core/n8450_6 ),
	.I2(\top/processor/sha_core/n8450_7 ),
	.I3(\top/processor/sha_core/n8450_8 ),
	.F(\top/processor/sha_core/n8450_4 )
);
defparam \top/processor/sha_core/n8450_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8451_s1  (
	.I0(\top/processor/sha_core/n8451_6 ),
	.I1(\top/processor/sha_core/n8451_7 ),
	.I2(\top/processor/sha_core/n8451_8 ),
	.I3(\top/processor/sha_core/n8451_9 ),
	.F(\top/processor/sha_core/n8451_4 )
);
defparam \top/processor/sha_core/n8451_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8451_s2  (
	.I0(\top/processor/sha_core/n8451_10 ),
	.I1(\top/processor/sha_core/n8451_11 ),
	.I2(\top/processor/sha_core/n8451_12 ),
	.I3(\top/processor/sha_core/n8451_13 ),
	.F(\top/processor/sha_core/n8451_5 )
);
defparam \top/processor/sha_core/n8451_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8452_s1  (
	.I0(\top/processor/sha_core/n8452_6 ),
	.I1(\top/processor/sha_core/n8452_7 ),
	.I2(\top/processor/sha_core/n8452_8 ),
	.I3(\top/processor/sha_core/n8452_9 ),
	.F(\top/processor/sha_core/n8452_4 )
);
defparam \top/processor/sha_core/n8452_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8452_s2  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [457]),
	.I2(\top/processor/sha_core/n8452_10 ),
	.I3(\top/processor/sha_core/n8452_11 ),
	.F(\top/processor/sha_core/n8452_5 )
);
defparam \top/processor/sha_core/n8452_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8453_s1  (
	.I0(\top/processor/sha_core/n8453_6 ),
	.I1(\top/processor/sha_core/n8453_7 ),
	.I2(\top/processor/sha_core/n8453_8 ),
	.I3(\top/processor/sha_core/n8453_9 ),
	.F(\top/processor/sha_core/n8453_4 )
);
defparam \top/processor/sha_core/n8453_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8453_s2  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [168]),
	.I2(\top/processor/sha_core/n8453_10 ),
	.I3(\top/processor/sha_core/n8453_11 ),
	.F(\top/processor/sha_core/n8453_5 )
);
defparam \top/processor/sha_core/n8453_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8454_s1  (
	.I0(\top/processor/sha_core/n8454_6 ),
	.I1(\top/processor/sha_core/n8454_7 ),
	.I2(\top/processor/sha_core/n8454_8 ),
	.I3(\top/processor/sha_core/n8454_9 ),
	.F(\top/processor/sha_core/n8454_4 )
);
defparam \top/processor/sha_core/n8454_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8454_s2  (
	.I0(\top/processor/sha_core/w[14]_31_9 ),
	.I1(\top/processor/core_block [39]),
	.I2(\top/processor/sha_core/n8454_10 ),
	.I3(\top/processor/sha_core/n8454_11 ),
	.F(\top/processor/sha_core/n8454_5 )
);
defparam \top/processor/sha_core/n8454_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8455_s1  (
	.I0(\top/processor/sha_core/n8455_6 ),
	.I1(\top/processor/sha_core/n8455_7 ),
	.I2(\top/processor/sha_core/n8455_8 ),
	.I3(\top/processor/sha_core/n8455_9 ),
	.F(\top/processor/sha_core/n8455_4 )
);
defparam \top/processor/sha_core/n8455_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8455_s2  (
	.I0(\top/processor/sha_core/n8455_10 ),
	.I1(\top/processor/sha_core/n8455_11 ),
	.I2(\top/processor/sha_core/n8455_12 ),
	.I3(\top/processor/sha_core/n8455_13 ),
	.F(\top/processor/sha_core/n8455_5 )
);
defparam \top/processor/sha_core/n8455_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8456_s1  (
	.I0(\top/processor/sha_core/n8456_6 ),
	.I1(\top/processor/sha_core/n8456_7 ),
	.I2(\top/processor/sha_core/n8456_8 ),
	.I3(\top/processor/sha_core/n8456_9 ),
	.F(\top/processor/sha_core/n8456_4 )
);
defparam \top/processor/sha_core/n8456_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8456_s2  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [261]),
	.I2(\top/processor/sha_core/n8456_10 ),
	.I3(\top/processor/sha_core/n8456_11 ),
	.F(\top/processor/sha_core/n8456_5 )
);
defparam \top/processor/sha_core/n8456_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8457_s1  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/core_block [228]),
	.I2(\top/processor/sha_core/n8457_5 ),
	.I3(\top/processor/sha_core/n8457_6 ),
	.F(\top/processor/sha_core/n8457_4 )
);
defparam \top/processor/sha_core/n8457_s1 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8458_s1  (
	.I0(\top/processor/sha_core/n8458_6 ),
	.I1(\top/processor/sha_core/n8458_7 ),
	.I2(\top/processor/sha_core/n8458_8 ),
	.I3(\top/processor/sha_core/n8458_9 ),
	.F(\top/processor/sha_core/n8458_4 )
);
defparam \top/processor/sha_core/n8458_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8458_s2  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [483]),
	.I2(\top/processor/sha_core/n8458_10 ),
	.I3(\top/processor/sha_core/n8458_11 ),
	.F(\top/processor/sha_core/n8458_5 )
);
defparam \top/processor/sha_core/n8458_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8459_s1  (
	.I0(\top/processor/sha_core/n8459_6 ),
	.I1(\top/processor/sha_core/n8459_7 ),
	.I2(\top/processor/sha_core/n8459_8 ),
	.I3(\top/processor/sha_core/n8459_9 ),
	.F(\top/processor/sha_core/n8459_4 )
);
defparam \top/processor/sha_core/n8459_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8459_s2  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [162]),
	.I2(\top/processor/sha_core/n8459_10 ),
	.I3(\top/processor/sha_core/n8459_11 ),
	.F(\top/processor/sha_core/n8459_5 )
);
defparam \top/processor/sha_core/n8459_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8460_s1  (
	.I0(\top/processor/sha_core/n8460_6 ),
	.I1(\top/processor/sha_core/n8460_7 ),
	.I2(\top/processor/sha_core/n8460_8 ),
	.I3(\top/processor/sha_core/n8460_9 ),
	.F(\top/processor/sha_core/n8460_4 )
);
defparam \top/processor/sha_core/n8460_s1 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8460_s2  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [129]),
	.I2(\top/processor/sha_core/n8460_10 ),
	.I3(\top/processor/sha_core/n8460_11 ),
	.F(\top/processor/sha_core/n8460_5 )
);
defparam \top/processor/sha_core/n8460_s2 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8461_s1  (
	.I0(\top/processor/sha_core/w[15]_31_11 ),
	.I1(\top/processor/core_block [0]),
	.I2(\top/processor/sha_core/n8461_6 ),
	.I3(\top/processor/sha_core/n8461_7 ),
	.F(\top/processor/sha_core/n8461_4 )
);
defparam \top/processor/sha_core/n8461_s1 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8461_s2  (
	.I0(\top/processor/sha_core/n8461_8 ),
	.I1(\top/processor/sha_core/n8461_9 ),
	.I2(\top/processor/sha_core/n8461_10 ),
	.I3(\top/processor/sha_core/n8461_11 ),
	.F(\top/processor/sha_core/n8461_5 )
);
defparam \top/processor/sha_core/n8461_s2 .INIT=16'h8000;
LUT3 \top/processor/sha_core/state_0_s4  (
	.I0(\top/processor/sha_core/t [6]),
	.I1(\top/processor/sha_core/msg_idx [6]),
	.I2(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/state_0_9 )
);
defparam \top/processor/sha_core/state_0_s4 .INIT=8'h3A;
LUT2 \top/processor/sha_core/w[0]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.F(\top/processor/sha_core/w[0]_31_9 )
);
defparam \top/processor/sha_core/w[0]_31_s5 .INIT=4'h1;
LUT4 \top/processor/sha_core/w[0]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[0]_31_10 )
);
defparam \top/processor/sha_core/w[0]_31_s6 .INIT=16'h0100;
LUT4 \top/processor/sha_core/w[1]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[1]_31_9 )
);
defparam \top/processor/sha_core/w[1]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[2]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [1]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/w[2]_31_9 )
);
defparam \top/processor/sha_core/w[2]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[3]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [1]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/w[3]_31_9 )
);
defparam \top/processor/sha_core/w[3]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[4]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/w[4]_31_9 )
);
defparam \top/processor/sha_core/w[4]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[5]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/w[5]_31_9 )
);
defparam \top/processor/sha_core/w[5]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[6]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/w[6]_31_9 )
);
defparam \top/processor/sha_core/w[6]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[8]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[8]_31_9 )
);
defparam \top/processor/sha_core/w[8]_31_s5 .INIT=16'h0100;
LUT4 \top/processor/sha_core/w[9]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[9]_31_9 )
);
defparam \top/processor/sha_core/w[9]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[10]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [1]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[10]_31_9 )
);
defparam \top/processor/sha_core/w[10]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[11]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [1]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[11]_31_9 )
);
defparam \top/processor/sha_core/w[11]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[12]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[12]_31_9 )
);
defparam \top/processor/sha_core/w[12]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[13]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[13]_31_9 )
);
defparam \top/processor/sha_core/w[13]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[14]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[14]_31_9 )
);
defparam \top/processor/sha_core/w[14]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[18]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [1]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[18]_31_9 )
);
defparam \top/processor/sha_core/w[18]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[19]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [2]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [1]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[19]_31_9 )
);
defparam \top/processor/sha_core/w[19]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[20]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[20]_31_9 )
);
defparam \top/processor/sha_core/w[20]_31_s5 .INIT=16'h1000;
LUT4 \top/processor/sha_core/w[21]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[21]_31_9 )
);
defparam \top/processor/sha_core/w[21]_31_s5 .INIT=16'h4000;
LUT4 \top/processor/sha_core/w[22]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [0]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[22]_31_9 )
);
defparam \top/processor/sha_core/w[22]_31_s5 .INIT=16'h4000;
LUT2 \top/processor/sha_core/w[40]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [3]),
	.F(\top/processor/sha_core/w[40]_31_9 )
);
defparam \top/processor/sha_core/w[40]_31_s5 .INIT=4'h4;
LUT3 \top/processor/sha_core/w[63]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [6]),
	.I1(\top/processor/sha_core/state [1]),
	.I2(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/w[63]_31_9 )
);
defparam \top/processor/sha_core/w[63]_31_s5 .INIT=8'h10;
LUT3 \top/processor/sha_core/n293_s5653  (
	.I0(\top/processor/sha_core/n293_7309 ),
	.I1(\top/processor/sha_core/n293_7310 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7225 )
);
defparam \top/processor/sha_core/n293_s5653 .INIT=8'h53;
LUT4 \top/processor/sha_core/n293_s5654  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/n293_7311 ),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7226 )
);
defparam \top/processor/sha_core/n293_s5654 .INIT=16'h35CB;
LUT4 \top/processor/sha_core/n293_s5655  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/n293_7312 ),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7227 )
);
defparam \top/processor/sha_core/n293_s5655 .INIT=16'h935C;
LUT3 \top/processor/sha_core/n293_s5656  (
	.I0(\top/processor/sha_core/n293_7313 ),
	.I1(\top/processor/sha_core/n293_7314 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7228 )
);
defparam \top/processor/sha_core/n293_s5656 .INIT=8'hC5;
LUT4 \top/processor/sha_core/n293_s5657  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7229 )
);
defparam \top/processor/sha_core/n293_s5657 .INIT=16'h4771;
LUT4 \top/processor/sha_core/n293_s5658  (
	.I0(\top/processor/sha_core/n293_7315 ),
	.I1(\top/processor/sha_core/n293_7316 ),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7230 )
);
defparam \top/processor/sha_core/n293_s5658 .INIT=16'hFA03;
LUT3 \top/processor/sha_core/n293_s5659  (
	.I0(\top/processor/sha_core/n293_7317 ),
	.I1(\top/processor/sha_core/t [0]),
	.I2(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7231 )
);
defparam \top/processor/sha_core/n293_s5659 .INIT=8'h10;
LUT4 \top/processor/sha_core/n293_s5660  (
	.I0(\top/processor/sha_core/n293_7318 ),
	.I1(\top/processor/sha_core/t [1]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7232 )
);
defparam \top/processor/sha_core/n293_s5660 .INIT=16'hE359;
LUT4 \top/processor/sha_core/n293_s5661  (
	.I0(\top/processor/sha_core/n293_7319 ),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/n293_7320 ),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7233 )
);
defparam \top/processor/sha_core/n293_s5661 .INIT=16'hBB0F;
LUT4 \top/processor/sha_core/n293_s5663  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7235 )
);
defparam \top/processor/sha_core/n293_s5663 .INIT=16'hE370;
LUT4 \top/processor/sha_core/n293_s5664  (
	.I0(\top/processor/sha_core/n293_7322 ),
	.I1(\top/processor/sha_core/n293_7388 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7236 )
);
defparam \top/processor/sha_core/n293_s5664 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n293_s5665  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/n293_7324 ),
	.F(\top/processor/sha_core/n293_7237 )
);
defparam \top/processor/sha_core/n293_s5665 .INIT=16'h5FC0;
LUT3 \top/processor/sha_core/n293_s5666  (
	.I0(\top/processor/sha_core/n293_7325 ),
	.I1(\top/processor/sha_core/n293_7326 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7238 )
);
defparam \top/processor/sha_core/n293_s5666 .INIT=8'hC5;
LUT4 \top/processor/sha_core/n293_s5667  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/n293_7327 ),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7239 )
);
defparam \top/processor/sha_core/n293_s5667 .INIT=16'hAC32;
LUT3 \top/processor/sha_core/n293_s5668  (
	.I0(\top/processor/sha_core/n293_7328 ),
	.I1(\top/processor/sha_core/n293_7329 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7240 )
);
defparam \top/processor/sha_core/n293_s5668 .INIT=8'hAC;
LUT4 \top/processor/sha_core/n293_s5669  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7241 )
);
defparam \top/processor/sha_core/n293_s5669 .INIT=16'h87FB;
LUT4 \top/processor/sha_core/n293_s5670  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7242 )
);
defparam \top/processor/sha_core/n293_s5670 .INIT=16'h68EE;
LUT4 \top/processor/sha_core/n293_s5671  (
	.I0(\top/processor/sha_core/n293_7330 ),
	.I1(\top/processor/sha_core/n293_7331 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7243 )
);
defparam \top/processor/sha_core/n293_s5671 .INIT=16'hF503;
LUT4 \top/processor/sha_core/n293_s5672  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7244 )
);
defparam \top/processor/sha_core/n293_s5672 .INIT=16'h419E;
LUT4 \top/processor/sha_core/n293_s5673  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7245 )
);
defparam \top/processor/sha_core/n293_s5673 .INIT=16'hBC44;
LUT4 \top/processor/sha_core/n293_s5674  (
	.I0(\top/processor/sha_core/n293_7332 ),
	.I1(\top/processor/sha_core/n293_7333 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7246 )
);
defparam \top/processor/sha_core/n293_s5674 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n293_s5675  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/n293_7334 ),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7247 )
);
defparam \top/processor/sha_core/n293_s5675 .INIT=16'hBC4B;
LUT4 \top/processor/sha_core/n293_s5676  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/n293_7335 ),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7248 )
);
defparam \top/processor/sha_core/n293_s5676 .INIT=16'h3D8F;
LUT4 \top/processor/sha_core/n293_s5677  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7249 )
);
defparam \top/processor/sha_core/n293_s5677 .INIT=16'hFC23;
LUT4 \top/processor/sha_core/n293_s5678  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7250 )
);
defparam \top/processor/sha_core/n293_s5678 .INIT=16'h4BB2;
LUT4 \top/processor/sha_core/n293_s5679  (
	.I0(\top/processor/sha_core/n293_7336 ),
	.I1(\top/processor/sha_core/n293_7337 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7251 )
);
defparam \top/processor/sha_core/n293_s5679 .INIT=16'h0CF5;
LUT4 \top/processor/sha_core/n293_s5680  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7252 )
);
defparam \top/processor/sha_core/n293_s5680 .INIT=16'h71EF;
LUT4 \top/processor/sha_core/n293_s5681  (
	.I0(\top/processor/sha_core/n293_7338 ),
	.I1(\top/processor/sha_core/n293_7339 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7253 )
);
defparam \top/processor/sha_core/n293_s5681 .INIT=16'h0CFA;
LUT4 \top/processor/sha_core/n293_s5682  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7254 )
);
defparam \top/processor/sha_core/n293_s5682 .INIT=16'hC5FB;
LUT4 \top/processor/sha_core/n293_s5683  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7255 )
);
defparam \top/processor/sha_core/n293_s5683 .INIT=16'h6BB0;
LUT4 \top/processor/sha_core/n293_s5684  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7256 )
);
defparam \top/processor/sha_core/n293_s5684 .INIT=16'hB5FC;
LUT4 \top/processor/sha_core/n293_s5685  (
	.I0(\top/processor/sha_core/n293_7340 ),
	.I1(\top/processor/sha_core/n293_7341 ),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7257 )
);
defparam \top/processor/sha_core/n293_s5685 .INIT=16'h0CF5;
LUT4 \top/processor/sha_core/n293_s5686  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7258 )
);
defparam \top/processor/sha_core/n293_s5686 .INIT=16'h310D;
LUT4 \top/processor/sha_core/n293_s5687  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7259 )
);
defparam \top/processor/sha_core/n293_s5687 .INIT=16'h30DF;
LUT4 \top/processor/sha_core/n293_s5688  (
	.I0(\top/processor/sha_core/n293_7342 ),
	.I1(\top/processor/sha_core/n293_7343 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7260 )
);
defparam \top/processor/sha_core/n293_s5688 .INIT=16'hF50C;
LUT4 \top/processor/sha_core/n293_s5689  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7261 )
);
defparam \top/processor/sha_core/n293_s5689 .INIT=16'h3CD4;
LUT4 \top/processor/sha_core/n293_s5690  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7262 )
);
defparam \top/processor/sha_core/n293_s5690 .INIT=16'h7F10;
LUT4 \top/processor/sha_core/n293_s5691  (
	.I0(\top/processor/sha_core/n293_7344 ),
	.I1(\top/processor/sha_core/n293_7345 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7263 )
);
defparam \top/processor/sha_core/n293_s5691 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n293_s5692  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7264 )
);
defparam \top/processor/sha_core/n293_s5692 .INIT=16'hCD5F;
LUT4 \top/processor/sha_core/n293_s5693  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7265 )
);
defparam \top/processor/sha_core/n293_s5693 .INIT=16'hF38E;
LUT4 \top/processor/sha_core/n293_s5694  (
	.I0(\top/processor/sha_core/n293_7346 ),
	.I1(\top/processor/sha_core/n293_7347 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7266 )
);
defparam \top/processor/sha_core/n293_s5694 .INIT=16'hF503;
LUT3 \top/processor/sha_core/n293_s5695  (
	.I0(\top/processor/sha_core/n293_7348 ),
	.I1(\top/processor/sha_core/n293_7349 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7267 )
);
defparam \top/processor/sha_core/n293_s5695 .INIT=8'h35;
LUT4 \top/processor/sha_core/n293_s5696  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/n293_7350 ),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7268 )
);
defparam \top/processor/sha_core/n293_s5696 .INIT=16'hC71E;
LUT4 \top/processor/sha_core/n293_s5697  (
	.I0(\top/processor/sha_core/n293_7351 ),
	.I1(\top/processor/sha_core/t [1]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7269 )
);
defparam \top/processor/sha_core/n293_s5697 .INIT=16'h94E8;
LUT3 \top/processor/sha_core/n293_s5698  (
	.I0(\top/processor/sha_core/n293_7352 ),
	.I1(\top/processor/sha_core/n293_7353 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7270 )
);
defparam \top/processor/sha_core/n293_s5698 .INIT=8'h53;
LUT4 \top/processor/sha_core/n293_s5699  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7271 )
);
defparam \top/processor/sha_core/n293_s5699 .INIT=16'h22CB;
LUT4 \top/processor/sha_core/n293_s5700  (
	.I0(\top/processor/sha_core/n293_7354 ),
	.I1(\top/processor/sha_core/n293_7355 ),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7272 )
);
defparam \top/processor/sha_core/n293_s5700 .INIT=16'h5FC0;
LUT4 \top/processor/sha_core/n293_s5701  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7273 )
);
defparam \top/processor/sha_core/n293_s5701 .INIT=16'hC3FA;
LUT4 \top/processor/sha_core/n293_s5702  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7274 )
);
defparam \top/processor/sha_core/n293_s5702 .INIT=16'hBE13;
LUT4 \top/processor/sha_core/n293_s5703  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7275 )
);
defparam \top/processor/sha_core/n293_s5703 .INIT=16'h4BFE;
LUT4 \top/processor/sha_core/n293_s5704  (
	.I0(\top/processor/sha_core/n293_7356 ),
	.I1(\top/processor/sha_core/n293_7357 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7276 )
);
defparam \top/processor/sha_core/n293_s5704 .INIT=16'h03F5;
LUT3 \top/processor/sha_core/n293_s5705  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7277 )
);
defparam \top/processor/sha_core/n293_s5705 .INIT=8'hD6;
LUT4 \top/processor/sha_core/n293_s5706  (
	.I0(\top/processor/sha_core/n293_7358 ),
	.I1(\top/processor/sha_core/n293_7359 ),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/t [0]),
	.F(\top/processor/sha_core/n293_7278 )
);
defparam \top/processor/sha_core/n293_s5706 .INIT=16'hAF30;
LUT4 \top/processor/sha_core/n293_s5707  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7279 )
);
defparam \top/processor/sha_core/n293_s5707 .INIT=16'hB6DF;
LUT4 \top/processor/sha_core/n293_s5708  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7280 )
);
defparam \top/processor/sha_core/n293_s5708 .INIT=16'h230E;
LUT4 \top/processor/sha_core/n293_s5709  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7281 )
);
defparam \top/processor/sha_core/n293_s5709 .INIT=16'h3F45;
LUT4 \top/processor/sha_core/n293_s5710  (
	.I0(\top/processor/sha_core/n293_7360 ),
	.I1(\top/processor/sha_core/n293_7361 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7282 )
);
defparam \top/processor/sha_core/n293_s5710 .INIT=16'h03F5;
LUT4 \top/processor/sha_core/n293_s5711  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7283 )
);
defparam \top/processor/sha_core/n293_s5711 .INIT=16'hD700;
LUT4 \top/processor/sha_core/n293_s5712  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7284 )
);
defparam \top/processor/sha_core/n293_s5712 .INIT=16'h9CA8;
LUT4 \top/processor/sha_core/n293_s5713  (
	.I0(\top/processor/sha_core/n293_7362 ),
	.I1(\top/processor/sha_core/n293_7363 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7285 )
);
defparam \top/processor/sha_core/n293_s5713 .INIT=16'h03F5;
LUT4 \top/processor/sha_core/n293_s5714  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/n293_7364 ),
	.F(\top/processor/sha_core/n293_7286 )
);
defparam \top/processor/sha_core/n293_s5714 .INIT=16'h007D;
LUT3 \top/processor/sha_core/n293_s5715  (
	.I0(\top/processor/sha_core/n293_7365 ),
	.I1(\top/processor/sha_core/n293_7366 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7287 )
);
defparam \top/processor/sha_core/n293_s5715 .INIT=8'h35;
LUT4 \top/processor/sha_core/n293_s5716  (
	.I0(\top/processor/sha_core/n293_7367 ),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7288 )
);
defparam \top/processor/sha_core/n293_s5716 .INIT=16'h2D8E;
LUT4 \top/processor/sha_core/n293_s5717  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/n293_7368 ),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7289 )
);
defparam \top/processor/sha_core/n293_s5717 .INIT=16'h038E;
LUT4 \top/processor/sha_core/n293_s5718  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7290 )
);
defparam \top/processor/sha_core/n293_s5718 .INIT=16'h789D;
LUT4 \top/processor/sha_core/n293_s5719  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7291 )
);
defparam \top/processor/sha_core/n293_s5719 .INIT=16'hDE03;
LUT4 \top/processor/sha_core/n293_s5720  (
	.I0(\top/processor/sha_core/n293_7369 ),
	.I1(\top/processor/sha_core/n293_7370 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7292 )
);
defparam \top/processor/sha_core/n293_s5720 .INIT=16'h03F5;
LUT4 \top/processor/sha_core/n293_s5721  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7293 )
);
defparam \top/processor/sha_core/n293_s5721 .INIT=16'hC4FC;
LUT4 \top/processor/sha_core/n293_s5722  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7294 )
);
defparam \top/processor/sha_core/n293_s5722 .INIT=16'hF832;
LUT4 \top/processor/sha_core/n293_s5723  (
	.I0(\top/processor/sha_core/n293_7371 ),
	.I1(\top/processor/sha_core/n293_7372 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7295 )
);
defparam \top/processor/sha_core/n293_s5723 .INIT=16'h0CF5;
LUT4 \top/processor/sha_core/n293_s5724  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7296 )
);
defparam \top/processor/sha_core/n293_s5724 .INIT=16'hA7FC;
LUT4 \top/processor/sha_core/n293_s5725  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7297 )
);
defparam \top/processor/sha_core/n293_s5725 .INIT=16'h45FC;
LUT4 \top/processor/sha_core/n293_s5726  (
	.I0(\top/processor/sha_core/n293_7373 ),
	.I1(\top/processor/sha_core/n293_7374 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7298 )
);
defparam \top/processor/sha_core/n293_s5726 .INIT=16'h03F5;
LUT3 \top/processor/sha_core/n293_s5727  (
	.I0(\top/processor/sha_core/n293_7375 ),
	.I1(\top/processor/sha_core/n293_7376 ),
	.I2(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7299 )
);
defparam \top/processor/sha_core/n293_s5727 .INIT=8'h5C;
LUT4 \top/processor/sha_core/n293_s5728  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/n293_7377 ),
	.F(\top/processor/sha_core/n293_7300 )
);
defparam \top/processor/sha_core/n293_s5728 .INIT=16'h0DF2;
LUT4 \top/processor/sha_core/n293_s5729  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/n293_7378 ),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7301 )
);
defparam \top/processor/sha_core/n293_s5729 .INIT=16'hE31E;
LUT4 \top/processor/sha_core/n293_s5730  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/n293_7379 ),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7302 )
);
defparam \top/processor/sha_core/n293_s5730 .INIT=16'hB2C3;
LUT4 \top/processor/sha_core/n293_s5731  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7303 )
);
defparam \top/processor/sha_core/n293_s5731 .INIT=16'hDD2F;
LUT4 \top/processor/sha_core/n293_s5732  (
	.I0(\top/processor/sha_core/n293_7380 ),
	.I1(\top/processor/sha_core/n293_7381 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7304 )
);
defparam \top/processor/sha_core/n293_s5732 .INIT=16'h30AF;
LUT4 \top/processor/sha_core/n293_s5733  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7305 )
);
defparam \top/processor/sha_core/n293_s5733 .INIT=16'h2C9B;
LUT4 \top/processor/sha_core/n293_s5734  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7306 )
);
defparam \top/processor/sha_core/n293_s5734 .INIT=16'h4F1B;
LUT4 \top/processor/sha_core/n293_s5735  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7307 )
);
defparam \top/processor/sha_core/n293_s5735 .INIT=16'hB645;
LUT4 \top/processor/sha_core/n293_s5736  (
	.I0(\top/processor/sha_core/n293_7382 ),
	.I1(\top/processor/sha_core/n293_7383 ),
	.I2(\top/processor/sha_core/t [0]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7308 )
);
defparam \top/processor/sha_core/n293_s5736 .INIT=16'hF50C;
LUT2 \top/processor/sha_core/n14441_s5  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/w[31]_31_11 ),
	.F(\top/processor/sha_core/n14441_10 )
);
defparam \top/processor/sha_core/n14441_s5 .INIT=4'h9;
LUT3 \top/processor/sha_core/n14439_s5  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/msg_idx [5]),
	.I2(\top/processor/sha_core/w[31]_31_11 ),
	.F(\top/processor/sha_core/n14439_10 )
);
defparam \top/processor/sha_core/n14439_s5 .INIT=8'h80;
LUT3 \top/processor/sha_core/n12131_s7  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [0]),
	.I2(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n12131_12 )
);
defparam \top/processor/sha_core/n12131_s7 .INIT=8'h80;
LUT3 \top/processor/sha_core/n12129_s7  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/n12131_12 ),
	.F(\top/processor/sha_core/n12129_12 )
);
defparam \top/processor/sha_core/n12129_s7 .INIT=8'h80;
LUT4 \top/processor/sha_core/n12128_s7  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/n12131_12 ),
	.F(\top/processor/sha_core/n12128_12 )
);
defparam \top/processor/sha_core/n12128_s7 .INIT=16'h8000;
LUT3 \top/processor/sha_core/n3578_s5  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.F(\top/processor/sha_core/n3578_12 )
);
defparam \top/processor/sha_core/n3578_s5 .INIT=8'h80;
LUT4 \top/processor/sha_core/n3766_s3  (
	.I0(\top/processor/sha_core/n3721_137 ),
	.I1(\top/processor/sha_core/n3721_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3766_11 ),
	.F(\top/processor/sha_core/n3766_6 )
);
defparam \top/processor/sha_core/n3766_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3766_s4  (
	.I0(\top/processor/sha_core/n3721_145 ),
	.I1(\top/processor/sha_core/n3721_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3766_12 ),
	.F(\top/processor/sha_core/n3766_7 )
);
defparam \top/processor/sha_core/n3766_s4 .INIT=16'hAFC0;
LUT3 \top/processor/sha_core/n3766_s5  (
	.I0(\top/processor/sha_core/msg_idx [4]),
	.I1(\top/processor/sha_core/w[31]_31_11 ),
	.I2(\top/processor/sha_core/msg_idx [5]),
	.F(\top/processor/sha_core/n3766_8 )
);
defparam \top/processor/sha_core/n3766_s5 .INIT=8'h1E;
LUT4 \top/processor/sha_core/n3766_s6  (
	.I0(\top/processor/sha_core/n3732_137 ),
	.I1(\top/processor/sha_core/n3732_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3766_13 ),
	.F(\top/processor/sha_core/n3766_9 )
);
defparam \top/processor/sha_core/n3766_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3766_s7  (
	.I0(\top/processor/sha_core/n3732_145 ),
	.I1(\top/processor/sha_core/n3732_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3766_14 ),
	.F(\top/processor/sha_core/n3766_10 )
);
defparam \top/processor/sha_core/n3766_s7 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3767_s3  (
	.I0(\top/processor/sha_core/n3720_137 ),
	.I1(\top/processor/sha_core/n3720_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3767_10 ),
	.F(\top/processor/sha_core/n3767_6 )
);
defparam \top/processor/sha_core/n3767_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3767_s4  (
	.I0(\top/processor/sha_core/n3720_145 ),
	.I1(\top/processor/sha_core/n3720_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3767_11 ),
	.F(\top/processor/sha_core/n3767_7 )
);
defparam \top/processor/sha_core/n3767_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3767_s5  (
	.I0(\top/processor/sha_core/n3731_137 ),
	.I1(\top/processor/sha_core/n3731_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3767_12 ),
	.F(\top/processor/sha_core/n3767_8 )
);
defparam \top/processor/sha_core/n3767_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3767_s6  (
	.I0(\top/processor/sha_core/n3731_145 ),
	.I1(\top/processor/sha_core/n3731_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3767_13 ),
	.F(\top/processor/sha_core/n3767_9 )
);
defparam \top/processor/sha_core/n3767_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3768_s3  (
	.I0(\top/processor/sha_core/n3719_137 ),
	.I1(\top/processor/sha_core/n3719_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3768_10 ),
	.F(\top/processor/sha_core/n3768_6 )
);
defparam \top/processor/sha_core/n3768_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3768_s4  (
	.I0(\top/processor/sha_core/n3719_145 ),
	.I1(\top/processor/sha_core/n3719_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3768_11 ),
	.F(\top/processor/sha_core/n3768_7 )
);
defparam \top/processor/sha_core/n3768_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3768_s5  (
	.I0(\top/processor/sha_core/n3730_137 ),
	.I1(\top/processor/sha_core/n3730_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3768_12 ),
	.F(\top/processor/sha_core/n3768_8 )
);
defparam \top/processor/sha_core/n3768_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3768_s6  (
	.I0(\top/processor/sha_core/n3730_145 ),
	.I1(\top/processor/sha_core/n3730_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3768_13 ),
	.F(\top/processor/sha_core/n3768_9 )
);
defparam \top/processor/sha_core/n3768_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3769_s4  (
	.I0(\top/processor/sha_core/n3718_137 ),
	.I1(\top/processor/sha_core/n3718_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3769_13 ),
	.F(\top/processor/sha_core/n3769_7 )
);
defparam \top/processor/sha_core/n3769_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3769_s5  (
	.I0(\top/processor/sha_core/n3718_145 ),
	.I1(\top/processor/sha_core/n3718_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3769_14 ),
	.F(\top/processor/sha_core/n3769_8 )
);
defparam \top/processor/sha_core/n3769_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3769_s6  (
	.I0(\top/processor/sha_core/n3729_137 ),
	.I1(\top/processor/sha_core/n3729_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3769_15 ),
	.F(\top/processor/sha_core/n3769_9 )
);
defparam \top/processor/sha_core/n3769_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3769_s7  (
	.I0(\top/processor/sha_core/n3729_145 ),
	.I1(\top/processor/sha_core/n3729_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3769_16 ),
	.F(\top/processor/sha_core/n3769_10 )
);
defparam \top/processor/sha_core/n3769_s7 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3769_s8  (
	.I0(\top/processor/sha_core/n3733_137 ),
	.I1(\top/processor/sha_core/n3733_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3769_17 ),
	.F(\top/processor/sha_core/n3769_11 )
);
defparam \top/processor/sha_core/n3769_s8 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3769_s9  (
	.I0(\top/processor/sha_core/n3733_145 ),
	.I1(\top/processor/sha_core/n3733_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3769_18 ),
	.F(\top/processor/sha_core/n3769_12 )
);
defparam \top/processor/sha_core/n3769_s9 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3770_s3  (
	.I0(\top/processor/sha_core/n3717_137 ),
	.I1(\top/processor/sha_core/n3717_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3770_10 ),
	.F(\top/processor/sha_core/n3770_6 )
);
defparam \top/processor/sha_core/n3770_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3770_s4  (
	.I0(\top/processor/sha_core/n3717_145 ),
	.I1(\top/processor/sha_core/n3717_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3770_11 ),
	.F(\top/processor/sha_core/n3770_7 )
);
defparam \top/processor/sha_core/n3770_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3770_s5  (
	.I0(\top/processor/sha_core/n3728_137 ),
	.I1(\top/processor/sha_core/n3728_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3770_12 ),
	.F(\top/processor/sha_core/n3770_8 )
);
defparam \top/processor/sha_core/n3770_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3770_s6  (
	.I0(\top/processor/sha_core/n3728_145 ),
	.I1(\top/processor/sha_core/n3728_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3770_13 ),
	.F(\top/processor/sha_core/n3770_9 )
);
defparam \top/processor/sha_core/n3770_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3771_s3  (
	.I0(\top/processor/sha_core/n3716_137 ),
	.I1(\top/processor/sha_core/n3716_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3771_10 ),
	.F(\top/processor/sha_core/n3771_6 )
);
defparam \top/processor/sha_core/n3771_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3771_s4  (
	.I0(\top/processor/sha_core/n3716_145 ),
	.I1(\top/processor/sha_core/n3716_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3771_11 ),
	.F(\top/processor/sha_core/n3771_7 )
);
defparam \top/processor/sha_core/n3771_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3771_s5  (
	.I0(\top/processor/sha_core/n3727_137 ),
	.I1(\top/processor/sha_core/n3727_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3771_12 ),
	.F(\top/processor/sha_core/n3771_8 )
);
defparam \top/processor/sha_core/n3771_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3771_s6  (
	.I0(\top/processor/sha_core/n3727_145 ),
	.I1(\top/processor/sha_core/n3727_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3771_13 ),
	.F(\top/processor/sha_core/n3771_9 )
);
defparam \top/processor/sha_core/n3771_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3772_s3  (
	.I0(\top/processor/sha_core/n3726_137 ),
	.I1(\top/processor/sha_core/n3726_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3772_10 ),
	.F(\top/processor/sha_core/n3772_6 )
);
defparam \top/processor/sha_core/n3772_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3772_s4  (
	.I0(\top/processor/sha_core/n3726_145 ),
	.I1(\top/processor/sha_core/n3726_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3772_11 ),
	.F(\top/processor/sha_core/n3772_7 )
);
defparam \top/processor/sha_core/n3772_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3772_s5  (
	.I0(\top/processor/sha_core/n3715_137 ),
	.I1(\top/processor/sha_core/n3715_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3772_12 ),
	.F(\top/processor/sha_core/n3772_8 )
);
defparam \top/processor/sha_core/n3772_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3772_s6  (
	.I0(\top/processor/sha_core/n3715_145 ),
	.I1(\top/processor/sha_core/n3715_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3772_13 ),
	.F(\top/processor/sha_core/n3772_9 )
);
defparam \top/processor/sha_core/n3772_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3773_s3  (
	.I0(\top/processor/sha_core/n3725_137 ),
	.I1(\top/processor/sha_core/n3725_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3773_10 ),
	.F(\top/processor/sha_core/n3773_6 )
);
defparam \top/processor/sha_core/n3773_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3773_s4  (
	.I0(\top/processor/sha_core/n3725_145 ),
	.I1(\top/processor/sha_core/n3725_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3773_11 ),
	.F(\top/processor/sha_core/n3773_7 )
);
defparam \top/processor/sha_core/n3773_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3773_s5  (
	.I0(\top/processor/sha_core/n3714_137 ),
	.I1(\top/processor/sha_core/n3714_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3773_12 ),
	.F(\top/processor/sha_core/n3773_8 )
);
defparam \top/processor/sha_core/n3773_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3773_s6  (
	.I0(\top/processor/sha_core/n3714_145 ),
	.I1(\top/processor/sha_core/n3714_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3773_13 ),
	.F(\top/processor/sha_core/n3773_9 )
);
defparam \top/processor/sha_core/n3773_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3774_s3  (
	.I0(\top/processor/sha_core/n3724_137 ),
	.I1(\top/processor/sha_core/n3724_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3774_10 ),
	.F(\top/processor/sha_core/n3774_6 )
);
defparam \top/processor/sha_core/n3774_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3774_s4  (
	.I0(\top/processor/sha_core/n3724_145 ),
	.I1(\top/processor/sha_core/n3724_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3774_11 ),
	.F(\top/processor/sha_core/n3774_7 )
);
defparam \top/processor/sha_core/n3774_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3774_s5  (
	.I0(\top/processor/sha_core/n3713_137 ),
	.I1(\top/processor/sha_core/n3713_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3774_12 ),
	.F(\top/processor/sha_core/n3774_8 )
);
defparam \top/processor/sha_core/n3774_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3774_s6  (
	.I0(\top/processor/sha_core/n3713_145 ),
	.I1(\top/processor/sha_core/n3713_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3774_13 ),
	.F(\top/processor/sha_core/n3774_9 )
);
defparam \top/processor/sha_core/n3774_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3775_s3  (
	.I0(\top/processor/sha_core/n3723_133 ),
	.I1(\top/processor/sha_core/n3723_137 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3775_10 ),
	.F(\top/processor/sha_core/n3775_6 )
);
defparam \top/processor/sha_core/n3775_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3775_s4  (
	.I0(\top/processor/sha_core/n3723_145 ),
	.I1(\top/processor/sha_core/n3723_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3775_11 ),
	.F(\top/processor/sha_core/n3775_7 )
);
defparam \top/processor/sha_core/n3775_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3775_s5  (
	.I0(\top/processor/sha_core/n3712_137 ),
	.I1(\top/processor/sha_core/n3712_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3775_12 ),
	.F(\top/processor/sha_core/n3775_8 )
);
defparam \top/processor/sha_core/n3775_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3775_s6  (
	.I0(\top/processor/sha_core/n3712_145 ),
	.I1(\top/processor/sha_core/n3712_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3775_13 ),
	.F(\top/processor/sha_core/n3775_9 )
);
defparam \top/processor/sha_core/n3775_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3776_s3  (
	.I0(\top/processor/sha_core/n3711_137 ),
	.I1(\top/processor/sha_core/n3711_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3776_10 ),
	.F(\top/processor/sha_core/n3776_6 )
);
defparam \top/processor/sha_core/n3776_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3776_s4  (
	.I0(\top/processor/sha_core/n3711_145 ),
	.I1(\top/processor/sha_core/n3711_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3776_11 ),
	.F(\top/processor/sha_core/n3776_7 )
);
defparam \top/processor/sha_core/n3776_s4 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3776_s5  (
	.I0(\top/processor/sha_core/n3722_137 ),
	.I1(\top/processor/sha_core/n3722_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3776_12 ),
	.F(\top/processor/sha_core/n3776_8 )
);
defparam \top/processor/sha_core/n3776_s5 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3776_s6  (
	.I0(\top/processor/sha_core/n3722_145 ),
	.I1(\top/processor/sha_core/n3722_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3776_13 ),
	.F(\top/processor/sha_core/n3776_9 )
);
defparam \top/processor/sha_core/n3776_s6 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3777_s2  (
	.I0(\top/processor/sha_core/n3710_137 ),
	.I1(\top/processor/sha_core/n3710_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3777_7 ),
	.F(\top/processor/sha_core/n3777_5 )
);
defparam \top/processor/sha_core/n3777_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3777_s3  (
	.I0(\top/processor/sha_core/n3710_145 ),
	.I1(\top/processor/sha_core/n3710_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3777_8 ),
	.F(\top/processor/sha_core/n3777_6 )
);
defparam \top/processor/sha_core/n3777_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3778_s2  (
	.I0(\top/processor/sha_core/n3709_137 ),
	.I1(\top/processor/sha_core/n3709_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3778_7 ),
	.F(\top/processor/sha_core/n3778_5 )
);
defparam \top/processor/sha_core/n3778_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3778_s3  (
	.I0(\top/processor/sha_core/n3709_145 ),
	.I1(\top/processor/sha_core/n3709_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3778_8 ),
	.F(\top/processor/sha_core/n3778_6 )
);
defparam \top/processor/sha_core/n3778_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3779_s2  (
	.I0(\top/processor/sha_core/n3708_137 ),
	.I1(\top/processor/sha_core/n3708_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3779_7 ),
	.F(\top/processor/sha_core/n3779_5 )
);
defparam \top/processor/sha_core/n3779_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3779_s3  (
	.I0(\top/processor/sha_core/n3708_145 ),
	.I1(\top/processor/sha_core/n3708_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3779_8 ),
	.F(\top/processor/sha_core/n3779_6 )
);
defparam \top/processor/sha_core/n3779_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3780_s2  (
	.I0(\top/processor/sha_core/n3707_137 ),
	.I1(\top/processor/sha_core/n3707_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3780_7 ),
	.F(\top/processor/sha_core/n3780_5 )
);
defparam \top/processor/sha_core/n3780_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3780_s3  (
	.I0(\top/processor/sha_core/n3707_145 ),
	.I1(\top/processor/sha_core/n3707_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3780_8 ),
	.F(\top/processor/sha_core/n3780_6 )
);
defparam \top/processor/sha_core/n3780_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3781_s2  (
	.I0(\top/processor/sha_core/n3706_137 ),
	.I1(\top/processor/sha_core/n3706_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3781_7 ),
	.F(\top/processor/sha_core/n3781_5 )
);
defparam \top/processor/sha_core/n3781_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3781_s3  (
	.I0(\top/processor/sha_core/n3706_145 ),
	.I1(\top/processor/sha_core/n3706_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3781_8 ),
	.F(\top/processor/sha_core/n3781_6 )
);
defparam \top/processor/sha_core/n3781_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3782_s2  (
	.I0(\top/processor/sha_core/n3705_137 ),
	.I1(\top/processor/sha_core/n3705_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3782_7 ),
	.F(\top/processor/sha_core/n3782_5 )
);
defparam \top/processor/sha_core/n3782_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3782_s3  (
	.I0(\top/processor/sha_core/n3705_145 ),
	.I1(\top/processor/sha_core/n3705_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3782_8 ),
	.F(\top/processor/sha_core/n3782_6 )
);
defparam \top/processor/sha_core/n3782_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3783_s2  (
	.I0(\top/processor/sha_core/n3736_137 ),
	.I1(\top/processor/sha_core/n3736_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3783_7 ),
	.F(\top/processor/sha_core/n3783_5 )
);
defparam \top/processor/sha_core/n3783_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3783_s3  (
	.I0(\top/processor/sha_core/n3736_145 ),
	.I1(\top/processor/sha_core/n3736_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3783_8 ),
	.F(\top/processor/sha_core/n3783_6 )
);
defparam \top/processor/sha_core/n3783_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3784_s2  (
	.I0(\top/processor/sha_core/n3735_137 ),
	.I1(\top/processor/sha_core/n3735_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3784_7 ),
	.F(\top/processor/sha_core/n3784_5 )
);
defparam \top/processor/sha_core/n3784_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3784_s3  (
	.I0(\top/processor/sha_core/n3735_145 ),
	.I1(\top/processor/sha_core/n3735_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3784_8 ),
	.F(\top/processor/sha_core/n3784_6 )
);
defparam \top/processor/sha_core/n3784_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3785_s2  (
	.I0(\top/processor/sha_core/n3734_137 ),
	.I1(\top/processor/sha_core/n3734_133 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3785_7 ),
	.F(\top/processor/sha_core/n3785_5 )
);
defparam \top/processor/sha_core/n3785_s2 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n3785_s3  (
	.I0(\top/processor/sha_core/n3734_145 ),
	.I1(\top/processor/sha_core/n3734_141 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n3785_8 ),
	.F(\top/processor/sha_core/n3785_6 )
);
defparam \top/processor/sha_core/n3785_s3 .INIT=16'hAFC0;
LUT4 \top/processor/sha_core/n8430_s4  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [287]),
	.I2(\top/processor/core_block [255]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8430_7 )
);
defparam \top/processor/sha_core/n8430_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8430_s5  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [351]),
	.I2(\top/processor/core_block [319]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8430_8 )
);
defparam \top/processor/sha_core/n8430_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8430_s6  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [223]),
	.I2(\top/processor/core_block [191]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8430_9 )
);
defparam \top/processor/sha_core/n8430_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8430_s7  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [159]),
	.I2(\top/processor/sha_core/n8430_14 ),
	.I3(\top/processor/sha_core/n8430_15 ),
	.F(\top/processor/sha_core/n8430_10 )
);
defparam \top/processor/sha_core/n8430_s7 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8430_s8  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/n8430_11 )
);
defparam \top/processor/sha_core/n8430_s8 .INIT=16'h0100;
LUT4 \top/processor/sha_core/n8430_s9  (
	.I0(\top/processor/core_block [415]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [383]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8430_12 )
);
defparam \top/processor/sha_core/n8430_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8430_s10  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [479]),
	.I2(\top/processor/core_block [447]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8430_13 )
);
defparam \top/processor/sha_core/n8430_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s3  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [2]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/n8431_6 )
);
defparam \top/processor/sha_core/n8431_s3 .INIT=16'h1000;
LUT4 \top/processor/sha_core/n8431_s4  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [510]),
	.I2(\top/processor/core_block [446]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8431_7 )
);
defparam \top/processor/sha_core/n8431_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s5  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [126]),
	.I2(\top/processor/sha_core/n8431_13 ),
	.I3(\top/processor/sha_core/n8431_14 ),
	.F(\top/processor/sha_core/n8431_8 )
);
defparam \top/processor/sha_core/n8431_s5 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8431_s6  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [222]),
	.I2(\top/processor/core_block [190]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8431_9 )
);
defparam \top/processor/sha_core/n8431_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s7  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [286]),
	.I2(\top/processor/core_block [254]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8431_10 )
);
defparam \top/processor/sha_core/n8431_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s8  (
	.I0(\top/processor/core_block [414]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [382]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8431_11 )
);
defparam \top/processor/sha_core/n8431_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s9  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [350]),
	.I2(\top/processor/core_block [318]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8431_12 )
);
defparam \top/processor/sha_core/n8431_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [349]),
	.I2(\top/processor/core_block [317]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8432_6 )
);
defparam \top/processor/sha_core/n8432_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s4  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [221]),
	.I2(\top/processor/core_block [189]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8432_7 )
);
defparam \top/processor/sha_core/n8432_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [285]),
	.I2(\top/processor/core_block [253]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8432_8 )
);
defparam \top/processor/sha_core/n8432_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [125]),
	.I2(\top/processor/sha_core/n8432_12 ),
	.I3(\top/processor/sha_core/n8432_13 ),
	.F(\top/processor/sha_core/n8432_9 )
);
defparam \top/processor/sha_core/n8432_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8432_s7  (
	.I0(\top/processor/core_block [445]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [381]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8432_10 )
);
defparam \top/processor/sha_core/n8432_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [509]),
	.I2(\top/processor/core_block [477]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8432_11 )
);
defparam \top/processor/sha_core/n8432_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [348]),
	.I2(\top/processor/core_block [316]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8433_6 )
);
defparam \top/processor/sha_core/n8433_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s4  (
	.I0(\top/processor/core_block [412]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [380]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8433_7 )
);
defparam \top/processor/sha_core/n8433_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [284]),
	.I2(\top/processor/core_block [252]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8433_8 )
);
defparam \top/processor/sha_core/n8433_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [124]),
	.I2(\top/processor/sha_core/n8433_12 ),
	.I3(\top/processor/sha_core/n8433_13 ),
	.F(\top/processor/sha_core/n8433_9 )
);
defparam \top/processor/sha_core/n8433_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8433_s7  (
	.I0(\top/processor/core_block [444]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [220]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8433_10 )
);
defparam \top/processor/sha_core/n8433_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [508]),
	.I2(\top/processor/core_block [476]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8433_11 )
);
defparam \top/processor/sha_core/n8433_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s3  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/core_block [251]),
	.I2(\top/processor/core_block [27]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8434_6 )
);
defparam \top/processor/sha_core/n8434_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [347]),
	.I2(\top/processor/core_block [59]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8434_7 )
);
defparam \top/processor/sha_core/n8434_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s5  (
	.I0(\top/processor/core_block [411]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [315]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8434_8 )
);
defparam \top/processor/sha_core/n8434_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s6  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [283]),
	.I2(\top/processor/core_block [91]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8434_9 )
);
defparam \top/processor/sha_core/n8434_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s7  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [219]),
	.I2(\top/processor/core_block [123]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8434_10 )
);
defparam \top/processor/sha_core/n8434_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [507]),
	.I2(\top/processor/sha_core/n8434_12 ),
	.I3(\top/processor/sha_core/n8434_13 ),
	.F(\top/processor/sha_core/n8434_11 )
);
defparam \top/processor/sha_core/n8434_s8 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8435_s3  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [90]),
	.I2(\top/processor/core_block [26]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8435_6 )
);
defparam \top/processor/sha_core/n8435_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s4  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [218]),
	.I2(\top/processor/core_block [122]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8435_7 )
);
defparam \top/processor/sha_core/n8435_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s5  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [154]),
	.I2(\top/processor/core_block [58]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8435_8 )
);
defparam \top/processor/sha_core/n8435_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s6  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [282]),
	.I2(\top/processor/core_block [186]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8435_9 )
);
defparam \top/processor/sha_core/n8435_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s7  (
	.I0(\top/processor/core_block [474]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [314]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8435_10 )
);
defparam \top/processor/sha_core/n8435_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s8  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [346]),
	.I2(\top/processor/core_block [250]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8435_11 )
);
defparam \top/processor/sha_core/n8435_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s9  (
	.I0(\top/processor/core_block [442]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [378]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8435_12 )
);
defparam \top/processor/sha_core/n8435_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8435_s10  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [506]),
	.I2(\top/processor/core_block [410]),
	.I3(\top/processor/sha_core/w[3]_31_9 ),
	.F(\top/processor/sha_core/n8435_13 )
);
defparam \top/processor/sha_core/n8435_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s3  (
	.I0(\top/processor/core_block [57]),
	.I1(\top/processor/sha_core/w[14]_31_9 ),
	.I2(\top/processor/core_block [25]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8436_6 )
);
defparam \top/processor/sha_core/n8436_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s4  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [281]),
	.I2(\top/processor/sha_core/n8436_12 ),
	.I3(\top/processor/sha_core/n8436_13 ),
	.F(\top/processor/sha_core/n8436_7 )
);
defparam \top/processor/sha_core/n8436_s4 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8436_s5  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [473]),
	.I2(\top/processor/core_block [441]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8436_8 )
);
defparam \top/processor/sha_core/n8436_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s6  (
	.I0(\top/processor/core_block [377]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [185]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8436_9 )
);
defparam \top/processor/sha_core/n8436_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s7  (
	.I0(\top/processor/core_block [505]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [217]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8436_10 )
);
defparam \top/processor/sha_core/n8436_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s8  (
	.I0(\top/processor/core_block [409]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [249]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8436_11 )
);
defparam \top/processor/sha_core/n8436_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [344]),
	.I2(\top/processor/core_block [312]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8437_6 )
);
defparam \top/processor/sha_core/n8437_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s4  (
	.I0(\top/processor/core_block [408]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [376]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8437_7 )
);
defparam \top/processor/sha_core/n8437_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [280]),
	.I2(\top/processor/core_block [248]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8437_8 )
);
defparam \top/processor/sha_core/n8437_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [120]),
	.I2(\top/processor/sha_core/n8437_12 ),
	.I3(\top/processor/sha_core/n8437_13 ),
	.F(\top/processor/sha_core/n8437_9 )
);
defparam \top/processor/sha_core/n8437_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8437_s7  (
	.I0(\top/processor/core_block [440]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [216]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8437_10 )
);
defparam \top/processor/sha_core/n8437_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [504]),
	.I2(\top/processor/core_block [472]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8437_11 )
);
defparam \top/processor/sha_core/n8437_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s3  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [311]),
	.I2(\top/processor/core_block [119]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8438_6 )
);
defparam \top/processor/sha_core/n8438_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s4  (
	.I0(\top/processor/core_block [407]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [343]),
	.I3(\top/processor/sha_core/w[5]_31_9 ),
	.F(\top/processor/sha_core/n8438_7 )
);
defparam \top/processor/sha_core/n8438_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s5  (
	.I0(\top/processor/core_block [439]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [215]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8438_8 )
);
defparam \top/processor/sha_core/n8438_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s6  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/core_block [247]),
	.I2(\top/processor/core_block [183]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8438_9 )
);
defparam \top/processor/sha_core/n8438_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s7  (
	.I0(\top/processor/core_block [375]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [23]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8438_10 )
);
defparam \top/processor/sha_core/n8438_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s8  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [151]),
	.I2(\top/processor/sha_core/n8438_12 ),
	.I3(\top/processor/sha_core/n8438_13 ),
	.F(\top/processor/sha_core/n8438_11 )
);
defparam \top/processor/sha_core/n8438_s8 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8439_s2  (
	.I0(\top/processor/sha_core/n8439_7 ),
	.I1(\top/processor/sha_core/n8439_8 ),
	.I2(\top/processor/sha_core/n8439_9 ),
	.I3(\top/processor/sha_core/n8439_10 ),
	.F(\top/processor/sha_core/n8439_5 )
);
defparam \top/processor/sha_core/n8439_s2 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8439_s3  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [310]),
	.I2(\top/processor/sha_core/n8439_11 ),
	.I3(\top/processor/sha_core/n8439_12 ),
	.F(\top/processor/sha_core/n8439_6 )
);
defparam \top/processor/sha_core/n8439_s3 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8440_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [341]),
	.I2(\top/processor/core_block [309]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8440_6 )
);
defparam \top/processor/sha_core/n8440_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8440_s4  (
	.I0(\top/processor/core_block [117]),
	.I1(\top/processor/sha_core/w[12]_31_9 ),
	.I2(\top/processor/core_block [21]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8440_7 )
);
defparam \top/processor/sha_core/n8440_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8440_s5  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [149]),
	.I2(\top/processor/core_block [53]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8440_8 )
);
defparam \top/processor/sha_core/n8440_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8440_s6  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [181]),
	.I2(\top/processor/sha_core/n8440_12 ),
	.I3(\top/processor/sha_core/n8440_13 ),
	.F(\top/processor/sha_core/n8440_9 )
);
defparam \top/processor/sha_core/n8440_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8440_s7  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [501]),
	.I2(\top/processor/core_block [469]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8440_10 )
);
defparam \top/processor/sha_core/n8440_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8440_s8  (
	.I0(\top/processor/core_block [437]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [373]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8440_11 )
);
defparam \top/processor/sha_core/n8440_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s3  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [276]),
	.I2(\top/processor/core_block [244]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8441_6 )
);
defparam \top/processor/sha_core/n8441_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [340]),
	.I2(\top/processor/core_block [308]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8441_7 )
);
defparam \top/processor/sha_core/n8441_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s5  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [212]),
	.I2(\top/processor/core_block [180]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8441_8 )
);
defparam \top/processor/sha_core/n8441_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [116]),
	.I2(\top/processor/sha_core/n8441_12 ),
	.I3(\top/processor/sha_core/n8441_13 ),
	.F(\top/processor/sha_core/n8441_9 )
);
defparam \top/processor/sha_core/n8441_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8441_s7  (
	.I0(\top/processor/core_block [404]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [372]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8441_10 )
);
defparam \top/processor/sha_core/n8441_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s8  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [468]),
	.I2(\top/processor/core_block [436]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8441_11 )
);
defparam \top/processor/sha_core/n8441_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8442_s2  (
	.I0(\top/processor/core_block [467]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [147]),
	.I3(\top/processor/sha_core/w[11]_31_9 ),
	.F(\top/processor/sha_core/n8442_5 )
);
defparam \top/processor/sha_core/n8442_s2 .INIT=16'h0777;
LUT3 \top/processor/sha_core/n8442_s3  (
	.I0(\top/processor/sha_core/w[14]_31_9 ),
	.I1(\top/processor/core_block [51]),
	.I2(\top/processor/sha_core/n8442_9 ),
	.F(\top/processor/sha_core/n8442_6 )
);
defparam \top/processor/sha_core/n8442_s3 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8442_s4  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/core_block [243]),
	.I2(\top/processor/sha_core/n8442_10 ),
	.I3(\top/processor/sha_core/n8442_11 ),
	.F(\top/processor/sha_core/n8442_7 )
);
defparam \top/processor/sha_core/n8442_s4 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8442_s5  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [83]),
	.I2(\top/processor/sha_core/n8442_12 ),
	.I3(\top/processor/sha_core/n8442_13 ),
	.F(\top/processor/sha_core/n8442_8 )
);
defparam \top/processor/sha_core/n8442_s5 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8443_s3  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [274]),
	.I2(\top/processor/core_block [242]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8443_6 )
);
defparam \top/processor/sha_core/n8443_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8443_s4  (
	.I0(\top/processor/core_block [402]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [18]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8443_7 )
);
defparam \top/processor/sha_core/n8443_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8443_s5  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [498]),
	.I2(\top/processor/core_block [466]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8443_8 )
);
defparam \top/processor/sha_core/n8443_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8443_s6  (
	.I0(\top/processor/sha_core/w[4]_31_9 ),
	.I1(\top/processor/core_block [370]),
	.I2(\top/processor/sha_core/n8443_12 ),
	.I3(\top/processor/sha_core/n8443_13 ),
	.F(\top/processor/sha_core/n8443_9 )
);
defparam \top/processor/sha_core/n8443_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8443_s7  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [338]),
	.I2(\top/processor/core_block [82]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8443_10 )
);
defparam \top/processor/sha_core/n8443_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8443_s8  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [210]),
	.I2(\top/processor/core_block [178]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8443_11 )
);
defparam \top/processor/sha_core/n8443_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s3  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [177]),
	.I2(\top/processor/core_block [17]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8444_6 )
);
defparam \top/processor/sha_core/n8444_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s4  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [273]),
	.I2(\top/processor/core_block [113]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8444_7 )
);
defparam \top/processor/sha_core/n8444_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s5  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [145]),
	.I2(\top/processor/core_block [49]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8444_8 )
);
defparam \top/processor/sha_core/n8444_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s6  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [209]),
	.I2(\top/processor/core_block [81]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8444_9 )
);
defparam \top/processor/sha_core/n8444_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s7  (
	.I0(\top/processor/core_block [433]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [305]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8444_10 )
);
defparam \top/processor/sha_core/n8444_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s8  (
	.I0(\top/processor/sha_core/w[4]_31_9 ),
	.I1(\top/processor/core_block [369]),
	.I2(\top/processor/sha_core/n8444_12 ),
	.I3(\top/processor/sha_core/n8444_13 ),
	.F(\top/processor/sha_core/n8444_11 )
);
defparam \top/processor/sha_core/n8444_s8 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8445_s3  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [496]),
	.I2(\top/processor/core_block [464]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8445_6 )
);
defparam \top/processor/sha_core/n8445_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s4  (
	.I0(\top/processor/core_block [400]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [336]),
	.I3(\top/processor/sha_core/w[5]_31_9 ),
	.F(\top/processor/sha_core/n8445_7 )
);
defparam \top/processor/sha_core/n8445_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s5  (
	.I0(\top/processor/core_block [432]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [368]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8445_8 )
);
defparam \top/processor/sha_core/n8445_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s6  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [304]),
	.I2(\top/processor/core_block [240]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8445_9 )
);
defparam \top/processor/sha_core/n8445_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s7  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [80]),
	.I2(\top/processor/core_block [16]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8445_10 )
);
defparam \top/processor/sha_core/n8445_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s8  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [208]),
	.I2(\top/processor/core_block [112]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8445_11 )
);
defparam \top/processor/sha_core/n8445_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [144]),
	.I2(\top/processor/core_block [48]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8445_12 )
);
defparam \top/processor/sha_core/n8445_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8445_s10  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [272]),
	.I2(\top/processor/core_block [176]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8445_13 )
);
defparam \top/processor/sha_core/n8445_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [335]),
	.I2(\top/processor/core_block [303]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8446_6 )
);
defparam \top/processor/sha_core/n8446_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s4  (
	.I0(\top/processor/core_block [399]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [367]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8446_7 )
);
defparam \top/processor/sha_core/n8446_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [271]),
	.I2(\top/processor/core_block [239]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8446_8 )
);
defparam \top/processor/sha_core/n8446_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s6  (
	.I0(\top/processor/sha_core/w[15]_31_11 ),
	.I1(\top/processor/core_block [15]),
	.I2(\top/processor/sha_core/n8446_12 ),
	.I3(\top/processor/sha_core/n8446_13 ),
	.F(\top/processor/sha_core/n8446_9 )
);
defparam \top/processor/sha_core/n8446_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8446_s7  (
	.I0(\top/processor/core_block [495]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [207]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8446_10 )
);
defparam \top/processor/sha_core/n8446_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s8  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [463]),
	.I2(\top/processor/core_block [431]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8446_11 )
);
defparam \top/processor/sha_core/n8446_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s3  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [462]),
	.I2(\top/processor/core_block [430]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8447_6 )
);
defparam \top/processor/sha_core/n8447_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s4  (
	.I0(\top/processor/core_block [366]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [14]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8447_7 )
);
defparam \top/processor/sha_core/n8447_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s5  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [78]),
	.I2(\top/processor/core_block [46]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8447_8 )
);
defparam \top/processor/sha_core/n8447_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s6  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [494]),
	.I2(\top/processor/sha_core/n8447_12 ),
	.I3(\top/processor/sha_core/n8447_13 ),
	.F(\top/processor/sha_core/n8447_9 )
);
defparam \top/processor/sha_core/n8447_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8447_s7  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [302]),
	.I2(\top/processor/core_block [174]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8447_10 )
);
defparam \top/processor/sha_core/n8447_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s8  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [270]),
	.I2(\top/processor/core_block [110]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8447_11 )
);
defparam \top/processor/sha_core/n8447_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s3  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [77]),
	.I2(\top/processor/core_block [13]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8448_6 )
);
defparam \top/processor/sha_core/n8448_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [333]),
	.I2(\top/processor/core_block [269]),
	.I3(\top/processor/sha_core/w[7]_31_11 ),
	.F(\top/processor/sha_core/n8448_7 )
);
defparam \top/processor/sha_core/n8448_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s5  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [301]),
	.I2(\top/processor/core_block [237]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8448_8 )
);
defparam \top/processor/sha_core/n8448_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s6  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [173]),
	.I2(\top/processor/sha_core/n8448_12 ),
	.I3(\top/processor/sha_core/n8448_13 ),
	.F(\top/processor/sha_core/n8448_9 )
);
defparam \top/processor/sha_core/n8448_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8448_s7  (
	.I0(\top/processor/core_block [461]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [365]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8448_10 )
);
defparam \top/processor/sha_core/n8448_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s8  (
	.I0(\top/processor/core_block [429]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [397]),
	.I3(\top/processor/sha_core/w[3]_31_9 ),
	.F(\top/processor/sha_core/n8448_11 )
);
defparam \top/processor/sha_core/n8448_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s3  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [268]),
	.I2(\top/processor/core_block [236]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8449_6 )
);
defparam \top/processor/sha_core/n8449_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [332]),
	.I2(\top/processor/core_block [204]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8449_7 )
);
defparam \top/processor/sha_core/n8449_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s5  (
	.I0(\top/processor/core_block [396]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [300]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8449_8 )
);
defparam \top/processor/sha_core/n8449_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s6  (
	.I0(\top/processor/core_block [428]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [108]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8449_9 )
);
defparam \top/processor/sha_core/n8449_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s7  (
	.I0(\top/processor/core_block [364]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [12]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8449_10 )
);
defparam \top/processor/sha_core/n8449_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s8  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [140]),
	.I2(\top/processor/sha_core/n8449_12 ),
	.I3(\top/processor/sha_core/n8449_13 ),
	.F(\top/processor/sha_core/n8449_11 )
);
defparam \top/processor/sha_core/n8449_s8 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8450_s2  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [267]),
	.I2(\top/processor/core_block [235]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8450_5 )
);
defparam \top/processor/sha_core/n8450_s2 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8450_s3  (
	.I0(\top/processor/sha_core/n8450_9 ),
	.I1(\top/processor/sha_core/n8450_10 ),
	.I2(\top/processor/sha_core/n8450_11 ),
	.I3(\top/processor/sha_core/n8450_12 ),
	.F(\top/processor/sha_core/n8450_6 )
);
defparam \top/processor/sha_core/n8450_s3 .INIT=16'h8000;
LUT3 \top/processor/sha_core/n8450_s4  (
	.I0(\top/processor/sha_core/w[3]_31_9 ),
	.I1(\top/processor/core_block [395]),
	.I2(\top/processor/sha_core/n8450_13 ),
	.F(\top/processor/sha_core/n8450_7 )
);
defparam \top/processor/sha_core/n8450_s4 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8450_s5  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [203]),
	.I2(\top/processor/core_block [171]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8450_8 )
);
defparam \top/processor/sha_core/n8450_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s3  (
	.I0(\top/processor/core_block [458]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [298]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8451_6 )
);
defparam \top/processor/sha_core/n8451_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [330]),
	.I2(\top/processor/core_block [234]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8451_7 )
);
defparam \top/processor/sha_core/n8451_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s5  (
	.I0(\top/processor/core_block [426]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [362]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8451_8 )
);
defparam \top/processor/sha_core/n8451_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s6  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [490]),
	.I2(\top/processor/core_block [394]),
	.I3(\top/processor/sha_core/w[3]_31_9 ),
	.F(\top/processor/sha_core/n8451_9 )
);
defparam \top/processor/sha_core/n8451_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s7  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [74]),
	.I2(\top/processor/core_block [10]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8451_10 )
);
defparam \top/processor/sha_core/n8451_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s8  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [202]),
	.I2(\top/processor/core_block [106]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8451_11 )
);
defparam \top/processor/sha_core/n8451_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [138]),
	.I2(\top/processor/core_block [42]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8451_12 )
);
defparam \top/processor/sha_core/n8451_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8451_s10  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [266]),
	.I2(\top/processor/core_block [170]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8451_13 )
);
defparam \top/processor/sha_core/n8451_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [329]),
	.I2(\top/processor/core_block [297]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8452_6 )
);
defparam \top/processor/sha_core/n8452_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s4  (
	.I0(\top/processor/core_block [393]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [361]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8452_7 )
);
defparam \top/processor/sha_core/n8452_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [265]),
	.I2(\top/processor/core_block [233]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8452_8 )
);
defparam \top/processor/sha_core/n8452_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [105]),
	.I2(\top/processor/sha_core/n8452_12 ),
	.I3(\top/processor/sha_core/n8452_13 ),
	.F(\top/processor/sha_core/n8452_9 )
);
defparam \top/processor/sha_core/n8452_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8452_s7  (
	.I0(\top/processor/core_block [425]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [169]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8452_10 )
);
defparam \top/processor/sha_core/n8452_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s8  (
	.I0(\top/processor/core_block [489]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [201]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8452_11 )
);
defparam \top/processor/sha_core/n8452_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [328]),
	.I2(\top/processor/core_block [296]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8453_6 )
);
defparam \top/processor/sha_core/n8453_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s4  (
	.I0(\top/processor/core_block [392]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [360]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8453_7 )
);
defparam \top/processor/sha_core/n8453_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [264]),
	.I2(\top/processor/core_block [232]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8453_8 )
);
defparam \top/processor/sha_core/n8453_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [104]),
	.I2(\top/processor/sha_core/n8453_12 ),
	.I3(\top/processor/sha_core/n8453_13 ),
	.F(\top/processor/sha_core/n8453_9 )
);
defparam \top/processor/sha_core/n8453_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8453_s7  (
	.I0(\top/processor/core_block [424]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [200]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8453_10 )
);
defparam \top/processor/sha_core/n8453_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [488]),
	.I2(\top/processor/core_block [456]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8453_11 )
);
defparam \top/processor/sha_core/n8453_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s3  (
	.I0(\top/processor/sha_core/w[8]_31_9 ),
	.I1(\top/processor/core_block [231]),
	.I2(\top/processor/core_block [103]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8454_6 )
);
defparam \top/processor/sha_core/n8454_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s4  (
	.I0(\top/processor/core_block [391]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [295]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8454_7 )
);
defparam \top/processor/sha_core/n8454_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s5  (
	.I0(\top/processor/core_block [423]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [199]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8454_8 )
);
defparam \top/processor/sha_core/n8454_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s6  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [327]),
	.I2(\top/processor/core_block [167]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8454_9 )
);
defparam \top/processor/sha_core/n8454_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s7  (
	.I0(\top/processor/core_block [359]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [7]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8454_10 )
);
defparam \top/processor/sha_core/n8454_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s8  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [135]),
	.I2(\top/processor/sha_core/n8454_12 ),
	.I3(\top/processor/sha_core/n8454_13 ),
	.F(\top/processor/sha_core/n8454_11 )
);
defparam \top/processor/sha_core/n8454_s8 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8455_s3  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [70]),
	.I2(\top/processor/core_block [6]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8455_6 )
);
defparam \top/processor/sha_core/n8455_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s4  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [198]),
	.I2(\top/processor/core_block [102]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8455_7 )
);
defparam \top/processor/sha_core/n8455_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s5  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [134]),
	.I2(\top/processor/core_block [38]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8455_8 )
);
defparam \top/processor/sha_core/n8455_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s6  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [262]),
	.I2(\top/processor/core_block [166]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8455_9 )
);
defparam \top/processor/sha_core/n8455_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s7  (
	.I0(\top/processor/core_block [454]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [358]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8455_10 )
);
defparam \top/processor/sha_core/n8455_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s8  (
	.I0(\top/processor/core_block [486]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [326]),
	.I3(\top/processor/sha_core/w[5]_31_9 ),
	.F(\top/processor/sha_core/n8455_11 )
);
defparam \top/processor/sha_core/n8455_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s9  (
	.I0(\top/processor/core_block [422]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [390]),
	.I3(\top/processor/sha_core/w[3]_31_9 ),
	.F(\top/processor/sha_core/n8455_12 )
);
defparam \top/processor/sha_core/n8455_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8455_s10  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [294]),
	.I2(\top/processor/core_block [230]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8455_13 )
);
defparam \top/processor/sha_core/n8455_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s3  (
	.I0(\top/processor/core_block [133]),
	.I1(\top/processor/sha_core/w[11]_31_9 ),
	.I2(\top/processor/core_block [69]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8456_6 )
);
defparam \top/processor/sha_core/n8456_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s4  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [293]),
	.I2(\top/processor/core_block [5]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8456_7 )
);
defparam \top/processor/sha_core/n8456_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s5  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [197]),
	.I2(\top/processor/core_block [101]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8456_8 )
);
defparam \top/processor/sha_core/n8456_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s6  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [165]),
	.I2(\top/processor/core_block [37]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8456_9 )
);
defparam \top/processor/sha_core/n8456_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s7  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [325]),
	.I2(\top/processor/core_block [229]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8456_10 )
);
defparam \top/processor/sha_core/n8456_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s8  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [453]),
	.I2(\top/processor/sha_core/n8456_12 ),
	.I3(\top/processor/sha_core/n8456_13 ),
	.F(\top/processor/sha_core/n8456_11 )
);
defparam \top/processor/sha_core/n8456_s8 .INIT=16'h7000;
LUT3 \top/processor/sha_core/n8457_s2  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [196]),
	.I2(\top/processor/sha_core/n8457_7 ),
	.F(\top/processor/sha_core/n8457_5 )
);
defparam \top/processor/sha_core/n8457_s2 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8457_s3  (
	.I0(\top/processor/sha_core/n8457_8 ),
	.I1(\top/processor/sha_core/n8457_9 ),
	.I2(\top/processor/sha_core/n8457_10 ),
	.I3(\top/processor/sha_core/n8457_11 ),
	.F(\top/processor/sha_core/n8457_6 )
);
defparam \top/processor/sha_core/n8457_s3 .INIT=16'h8000;
LUT4 \top/processor/sha_core/n8458_s3  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [259]),
	.I2(\top/processor/core_block [227]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8458_6 )
);
defparam \top/processor/sha_core/n8458_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8458_s4  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [323]),
	.I2(\top/processor/core_block [291]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8458_7 )
);
defparam \top/processor/sha_core/n8458_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8458_s5  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [195]),
	.I2(\top/processor/core_block [163]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8458_8 )
);
defparam \top/processor/sha_core/n8458_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8458_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [99]),
	.I2(\top/processor/sha_core/n8458_12 ),
	.I3(\top/processor/sha_core/n8458_13 ),
	.F(\top/processor/sha_core/n8458_9 )
);
defparam \top/processor/sha_core/n8458_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8458_s7  (
	.I0(\top/processor/core_block [387]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [355]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8458_10 )
);
defparam \top/processor/sha_core/n8458_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8458_s8  (
	.I0(\top/processor/sha_core/n8431_6 ),
	.I1(\top/processor/core_block [451]),
	.I2(\top/processor/core_block [419]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8458_11 )
);
defparam \top/processor/sha_core/n8458_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s3  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [322]),
	.I2(\top/processor/core_block [290]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8459_6 )
);
defparam \top/processor/sha_core/n8459_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s4  (
	.I0(\top/processor/core_block [386]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [354]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8459_7 )
);
defparam \top/processor/sha_core/n8459_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s5  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [258]),
	.I2(\top/processor/core_block [226]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8459_8 )
);
defparam \top/processor/sha_core/n8459_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s6  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [98]),
	.I2(\top/processor/sha_core/n8459_12 ),
	.I3(\top/processor/sha_core/n8459_13 ),
	.F(\top/processor/sha_core/n8459_9 )
);
defparam \top/processor/sha_core/n8459_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8459_s7  (
	.I0(\top/processor/core_block [418]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [194]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8459_10 )
);
defparam \top/processor/sha_core/n8459_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [482]),
	.I2(\top/processor/core_block [450]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8459_11 )
);
defparam \top/processor/sha_core/n8459_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s3  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [289]),
	.I2(\top/processor/core_block [225]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8460_6 )
);
defparam \top/processor/sha_core/n8460_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s4  (
	.I0(\top/processor/core_block [481]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [321]),
	.I3(\top/processor/sha_core/w[5]_31_9 ),
	.F(\top/processor/sha_core/n8460_7 )
);
defparam \top/processor/sha_core/n8460_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s5  (
	.I0(\top/processor/core_block [449]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [65]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8460_8 )
);
defparam \top/processor/sha_core/n8460_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s6  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [161]),
	.I2(\top/processor/sha_core/n8460_12 ),
	.I3(\top/processor/sha_core/n8460_13 ),
	.F(\top/processor/sha_core/n8460_9 )
);
defparam \top/processor/sha_core/n8460_s6 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8460_s7  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [257]),
	.I2(\top/processor/core_block [1]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8460_10 )
);
defparam \top/processor/sha_core/n8460_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s8  (
	.I0(\top/processor/core_block [353]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [33]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8460_11 )
);
defparam \top/processor/sha_core/n8460_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s3  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [128]),
	.I2(\top/processor/core_block [32]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8461_6 )
);
defparam \top/processor/sha_core/n8461_s3 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s4  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [64]),
	.I2(\top/processor/sha_core/n8461_12 ),
	.I3(\top/processor/sha_core/n8461_13 ),
	.F(\top/processor/sha_core/n8461_7 )
);
defparam \top/processor/sha_core/n8461_s4 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8461_s5  (
	.I0(\top/processor/core_block [384]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [288]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8461_8 )
);
defparam \top/processor/sha_core/n8461_s5 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s6  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [480]),
	.I2(\top/processor/core_block [416]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8461_9 )
);
defparam \top/processor/sha_core/n8461_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s7  (
	.I0(\top/processor/core_block [448]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [352]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8461_10 )
);
defparam \top/processor/sha_core/n8461_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s8  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [320]),
	.I2(\top/processor/core_block [224]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8461_11 )
);
defparam \top/processor/sha_core/n8461_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n293_s5737  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7309 )
);
defparam \top/processor/sha_core/n293_s5737 .INIT=16'h15FE;
LUT4 \top/processor/sha_core/n293_s5738  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7310 )
);
defparam \top/processor/sha_core/n293_s5738 .INIT=16'hB42B;
LUT3 \top/processor/sha_core/n293_s5739  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [1]),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7311 )
);
defparam \top/processor/sha_core/n293_s5739 .INIT=8'h90;
LUT4 \top/processor/sha_core/n293_s5740  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7312 )
);
defparam \top/processor/sha_core/n293_s5740 .INIT=16'h1A47;
LUT4 \top/processor/sha_core/n293_s5741  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7313 )
);
defparam \top/processor/sha_core/n293_s5741 .INIT=16'hBCCA;
LUT4 \top/processor/sha_core/n293_s5742  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7314 )
);
defparam \top/processor/sha_core/n293_s5742 .INIT=16'h33C5;
LUT4 \top/processor/sha_core/n293_s5743  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7315 )
);
defparam \top/processor/sha_core/n293_s5743 .INIT=16'h71C0;
LUT4 \top/processor/sha_core/n293_s5744  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7316 )
);
defparam \top/processor/sha_core/n293_s5744 .INIT=16'hCBA7;
LUT3 \top/processor/sha_core/n293_s5745  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7317 )
);
defparam \top/processor/sha_core/n293_s5745 .INIT=8'hE3;
LUT4 \top/processor/sha_core/n293_s5746  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7318 )
);
defparam \top/processor/sha_core/n293_s5746 .INIT=16'h15E3;
LUT3 \top/processor/sha_core/n293_s5747  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7319 )
);
defparam \top/processor/sha_core/n293_s5747 .INIT=8'hBC;
LUT4 \top/processor/sha_core/n293_s5748  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7320 )
);
defparam \top/processor/sha_core/n293_s5748 .INIT=16'hBF68;
LUT4 \top/processor/sha_core/n293_s5750  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7322 )
);
defparam \top/processor/sha_core/n293_s5750 .INIT=16'hAC32;
LUT4 \top/processor/sha_core/n293_s5752  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7324 )
);
defparam \top/processor/sha_core/n293_s5752 .INIT=16'h2EE8;
LUT4 \top/processor/sha_core/n293_s5753  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7325 )
);
defparam \top/processor/sha_core/n293_s5753 .INIT=16'hBC4E;
LUT4 \top/processor/sha_core/n293_s5754  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7326 )
);
defparam \top/processor/sha_core/n293_s5754 .INIT=16'h453E;
LUT4 \top/processor/sha_core/n293_s5755  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7327 )
);
defparam \top/processor/sha_core/n293_s5755 .INIT=16'h2CEA;
LUT4 \top/processor/sha_core/n293_s5756  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7328 )
);
defparam \top/processor/sha_core/n293_s5756 .INIT=16'hA8FE;
LUT4 \top/processor/sha_core/n293_s5757  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7329 )
);
defparam \top/processor/sha_core/n293_s5757 .INIT=16'hEA2C;
LUT4 \top/processor/sha_core/n293_s5758  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7330 )
);
defparam \top/processor/sha_core/n293_s5758 .INIT=16'hC71F;
LUT4 \top/processor/sha_core/n293_s5759  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7331 )
);
defparam \top/processor/sha_core/n293_s5759 .INIT=16'hE09F;
LUT4 \top/processor/sha_core/n293_s5760  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7332 )
);
defparam \top/processor/sha_core/n293_s5760 .INIT=16'h9FF3;
LUT4 \top/processor/sha_core/n293_s5761  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7333 )
);
defparam \top/processor/sha_core/n293_s5761 .INIT=16'hB24B;
LUT4 \top/processor/sha_core/n293_s5762  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [1]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7334 )
);
defparam \top/processor/sha_core/n293_s5762 .INIT=16'hEC30;
LUT4 \top/processor/sha_core/n293_s5763  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [1]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7335 )
);
defparam \top/processor/sha_core/n293_s5763 .INIT=16'h453C;
LUT4 \top/processor/sha_core/n293_s5764  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7336 )
);
defparam \top/processor/sha_core/n293_s5764 .INIT=16'h4BFE;
LUT4 \top/processor/sha_core/n293_s5765  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7337 )
);
defparam \top/processor/sha_core/n293_s5765 .INIT=16'h1B54;
LUT4 \top/processor/sha_core/n293_s5766  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7338 )
);
defparam \top/processor/sha_core/n293_s5766 .INIT=16'hF1CF;
LUT4 \top/processor/sha_core/n293_s5767  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7339 )
);
defparam \top/processor/sha_core/n293_s5767 .INIT=16'h3D23;
LUT4 \top/processor/sha_core/n293_s5768  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7340 )
);
defparam \top/processor/sha_core/n293_s5768 .INIT=16'h6BF7;
LUT4 \top/processor/sha_core/n293_s5769  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7341 )
);
defparam \top/processor/sha_core/n293_s5769 .INIT=16'h00B2;
LUT4 \top/processor/sha_core/n293_s5770  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7342 )
);
defparam \top/processor/sha_core/n293_s5770 .INIT=16'hD8E3;
LUT4 \top/processor/sha_core/n293_s5771  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7343 )
);
defparam \top/processor/sha_core/n293_s5771 .INIT=16'h71CA;
LUT4 \top/processor/sha_core/n293_s5772  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7344 )
);
defparam \top/processor/sha_core/n293_s5772 .INIT=16'h95DC;
LUT4 \top/processor/sha_core/n293_s5773  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7345 )
);
defparam \top/processor/sha_core/n293_s5773 .INIT=16'h7807;
LUT4 \top/processor/sha_core/n293_s5774  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7346 )
);
defparam \top/processor/sha_core/n293_s5774 .INIT=16'h74A4;
LUT4 \top/processor/sha_core/n293_s5775  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7347 )
);
defparam \top/processor/sha_core/n293_s5775 .INIT=16'h7635;
LUT4 \top/processor/sha_core/n293_s5776  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7348 )
);
defparam \top/processor/sha_core/n293_s5776 .INIT=16'hBCAB;
LUT4 \top/processor/sha_core/n293_s5777  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7349 )
);
defparam \top/processor/sha_core/n293_s5777 .INIT=16'h7EC5;
LUT4 \top/processor/sha_core/n293_s5778  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [1]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7350 )
);
defparam \top/processor/sha_core/n293_s5778 .INIT=16'hDE3D;
LUT4 \top/processor/sha_core/n293_s5779  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7351 )
);
defparam \top/processor/sha_core/n293_s5779 .INIT=16'hCD5E;
LUT4 \top/processor/sha_core/n293_s5780  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7352 )
);
defparam \top/processor/sha_core/n293_s5780 .INIT=16'hA73F;
LUT4 \top/processor/sha_core/n293_s5781  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7353 )
);
defparam \top/processor/sha_core/n293_s5781 .INIT=16'hCBA0;
LUT4 \top/processor/sha_core/n293_s5782  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7354 )
);
defparam \top/processor/sha_core/n293_s5782 .INIT=16'h2C17;
LUT4 \top/processor/sha_core/n293_s5783  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7355 )
);
defparam \top/processor/sha_core/n293_s5783 .INIT=16'hB4FB;
LUT4 \top/processor/sha_core/n293_s5784  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7356 )
);
defparam \top/processor/sha_core/n293_s5784 .INIT=16'h9EE3;
LUT4 \top/processor/sha_core/n293_s5785  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7357 )
);
defparam \top/processor/sha_core/n293_s5785 .INIT=16'hEFB0;
LUT4 \top/processor/sha_core/n293_s5786  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7358 )
);
defparam \top/processor/sha_core/n293_s5786 .INIT=16'h6B90;
LUT4 \top/processor/sha_core/n293_s5787  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7359 )
);
defparam \top/processor/sha_core/n293_s5787 .INIT=16'h883A;
LUT4 \top/processor/sha_core/n293_s5788  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7360 )
);
defparam \top/processor/sha_core/n293_s5788 .INIT=16'h7817;
LUT4 \top/processor/sha_core/n293_s5789  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7361 )
);
defparam \top/processor/sha_core/n293_s5789 .INIT=16'h7EE3;
LUT4 \top/processor/sha_core/n293_s5790  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7362 )
);
defparam \top/processor/sha_core/n293_s5790 .INIT=16'h0B00;
LUT4 \top/processor/sha_core/n293_s5791  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7363 )
);
defparam \top/processor/sha_core/n293_s5791 .INIT=16'hBC4B;
LUT4 \top/processor/sha_core/n293_s5792  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7364 )
);
defparam \top/processor/sha_core/n293_s5792 .INIT=16'h6C53;
LUT4 \top/processor/sha_core/n293_s5793  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7365 )
);
defparam \top/processor/sha_core/n293_s5793 .INIT=16'h9671;
LUT4 \top/processor/sha_core/n293_s5794  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7366 )
);
defparam \top/processor/sha_core/n293_s5794 .INIT=16'hED3E;
LUT3 \top/processor/sha_core/n293_s5795  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7367 )
);
defparam \top/processor/sha_core/n293_s5795 .INIT=8'h70;
LUT4 \top/processor/sha_core/n293_s5796  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [1]),
	.F(\top/processor/sha_core/n293_7368 )
);
defparam \top/processor/sha_core/n293_s5796 .INIT=16'hB563;
LUT4 \top/processor/sha_core/n293_s5797  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7369 )
);
defparam \top/processor/sha_core/n293_s5797 .INIT=16'hF5CE;
LUT4 \top/processor/sha_core/n293_s5798  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7370 )
);
defparam \top/processor/sha_core/n293_s5798 .INIT=16'h349B;
LUT4 \top/processor/sha_core/n293_s5799  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7371 )
);
defparam \top/processor/sha_core/n293_s5799 .INIT=16'hBC4F;
LUT4 \top/processor/sha_core/n293_s5800  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7372 )
);
defparam \top/processor/sha_core/n293_s5800 .INIT=16'hCBA7;
LUT4 \top/processor/sha_core/n293_s5801  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7373 )
);
defparam \top/processor/sha_core/n293_s5801 .INIT=16'hF5C3;
LUT4 \top/processor/sha_core/n293_s5802  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7374 )
);
defparam \top/processor/sha_core/n293_s5802 .INIT=16'h5EC7;
LUT4 \top/processor/sha_core/n293_s5803  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7375 )
);
defparam \top/processor/sha_core/n293_s5803 .INIT=16'h9CC5;
LUT4 \top/processor/sha_core/n293_s5804  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7376 )
);
defparam \top/processor/sha_core/n293_s5804 .INIT=16'h07D1;
LUT4 \top/processor/sha_core/n293_s5805  (
	.I0(\top/processor/sha_core/t [1]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7377 )
);
defparam \top/processor/sha_core/n293_s5805 .INIT=16'h07E8;
LUT4 \top/processor/sha_core/n293_s5806  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [4]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [2]),
	.F(\top/processor/sha_core/n293_7378 )
);
defparam \top/processor/sha_core/n293_s5806 .INIT=16'h1FF3;
LUT4 \top/processor/sha_core/n293_s5807  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7379 )
);
defparam \top/processor/sha_core/n293_s5807 .INIT=16'h620B;
LUT4 \top/processor/sha_core/n293_s5808  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [3]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7380 )
);
defparam \top/processor/sha_core/n293_s5808 .INIT=16'h9370;
LUT4 \top/processor/sha_core/n293_s5809  (
	.I0(\top/processor/sha_core/t [5]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7381 )
);
defparam \top/processor/sha_core/n293_s5809 .INIT=16'hB04F;
LUT4 \top/processor/sha_core/n293_s5810  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [2]),
	.I2(\top/processor/sha_core/t [5]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7382 )
);
defparam \top/processor/sha_core/n293_s5810 .INIT=16'h09BA;
LUT4 \top/processor/sha_core/n293_s5811  (
	.I0(\top/processor/sha_core/t [3]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [4]),
	.F(\top/processor/sha_core/n293_7383 )
);
defparam \top/processor/sha_core/n293_s5811 .INIT=16'hA38A;
LUT4 \top/processor/sha_core/n3766_s8  (
	.I0(\top/processor/sha_core/n3721_139 ),
	.I1(\top/processor/sha_core/n3721_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3766_11 )
);
defparam \top/processor/sha_core/n3766_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3766_s9  (
	.I0(\top/processor/sha_core/n3721_147 ),
	.I1(\top/processor/sha_core/n3721_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3766_12 )
);
defparam \top/processor/sha_core/n3766_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3766_s10  (
	.I0(\top/processor/sha_core/n3732_139 ),
	.I1(\top/processor/sha_core/n3732_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3766_13 )
);
defparam \top/processor/sha_core/n3766_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3766_s11  (
	.I0(\top/processor/sha_core/n3732_147 ),
	.I1(\top/processor/sha_core/n3732_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3766_14 )
);
defparam \top/processor/sha_core/n3766_s11 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3767_s7  (
	.I0(\top/processor/sha_core/n3720_139 ),
	.I1(\top/processor/sha_core/n3720_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3767_10 )
);
defparam \top/processor/sha_core/n3767_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3767_s8  (
	.I0(\top/processor/sha_core/n3720_147 ),
	.I1(\top/processor/sha_core/n3720_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3767_11 )
);
defparam \top/processor/sha_core/n3767_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3767_s9  (
	.I0(\top/processor/sha_core/n3731_139 ),
	.I1(\top/processor/sha_core/n3731_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3767_12 )
);
defparam \top/processor/sha_core/n3767_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3767_s10  (
	.I0(\top/processor/sha_core/n3731_147 ),
	.I1(\top/processor/sha_core/n3731_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3767_13 )
);
defparam \top/processor/sha_core/n3767_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3768_s7  (
	.I0(\top/processor/sha_core/n3719_139 ),
	.I1(\top/processor/sha_core/n3719_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3768_10 )
);
defparam \top/processor/sha_core/n3768_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3768_s8  (
	.I0(\top/processor/sha_core/n3719_147 ),
	.I1(\top/processor/sha_core/n3719_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3768_11 )
);
defparam \top/processor/sha_core/n3768_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3768_s9  (
	.I0(\top/processor/sha_core/n3730_139 ),
	.I1(\top/processor/sha_core/n3730_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3768_12 )
);
defparam \top/processor/sha_core/n3768_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3768_s10  (
	.I0(\top/processor/sha_core/n3730_147 ),
	.I1(\top/processor/sha_core/n3730_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3768_13 )
);
defparam \top/processor/sha_core/n3768_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3769_s10  (
	.I0(\top/processor/sha_core/n3718_139 ),
	.I1(\top/processor/sha_core/n3718_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3769_13 )
);
defparam \top/processor/sha_core/n3769_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3769_s11  (
	.I0(\top/processor/sha_core/n3718_147 ),
	.I1(\top/processor/sha_core/n3718_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3769_14 )
);
defparam \top/processor/sha_core/n3769_s11 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3769_s12  (
	.I0(\top/processor/sha_core/n3729_139 ),
	.I1(\top/processor/sha_core/n3729_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3769_15 )
);
defparam \top/processor/sha_core/n3769_s12 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3769_s13  (
	.I0(\top/processor/sha_core/n3729_147 ),
	.I1(\top/processor/sha_core/n3729_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3769_16 )
);
defparam \top/processor/sha_core/n3769_s13 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3769_s14  (
	.I0(\top/processor/sha_core/n3733_139 ),
	.I1(\top/processor/sha_core/n3733_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3769_17 )
);
defparam \top/processor/sha_core/n3769_s14 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3769_s15  (
	.I0(\top/processor/sha_core/n3733_147 ),
	.I1(\top/processor/sha_core/n3733_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3769_18 )
);
defparam \top/processor/sha_core/n3769_s15 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3770_s7  (
	.I0(\top/processor/sha_core/n3717_139 ),
	.I1(\top/processor/sha_core/n3717_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3770_10 )
);
defparam \top/processor/sha_core/n3770_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3770_s8  (
	.I0(\top/processor/sha_core/n3717_147 ),
	.I1(\top/processor/sha_core/n3717_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3770_11 )
);
defparam \top/processor/sha_core/n3770_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3770_s9  (
	.I0(\top/processor/sha_core/n3728_139 ),
	.I1(\top/processor/sha_core/n3728_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3770_12 )
);
defparam \top/processor/sha_core/n3770_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3770_s10  (
	.I0(\top/processor/sha_core/n3728_147 ),
	.I1(\top/processor/sha_core/n3728_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3770_13 )
);
defparam \top/processor/sha_core/n3770_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3771_s7  (
	.I0(\top/processor/sha_core/n3716_139 ),
	.I1(\top/processor/sha_core/n3716_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3771_10 )
);
defparam \top/processor/sha_core/n3771_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3771_s8  (
	.I0(\top/processor/sha_core/n3716_147 ),
	.I1(\top/processor/sha_core/n3716_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3771_11 )
);
defparam \top/processor/sha_core/n3771_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3771_s9  (
	.I0(\top/processor/sha_core/n3727_139 ),
	.I1(\top/processor/sha_core/n3727_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3771_12 )
);
defparam \top/processor/sha_core/n3771_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3771_s10  (
	.I0(\top/processor/sha_core/n3727_147 ),
	.I1(\top/processor/sha_core/n3727_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3771_13 )
);
defparam \top/processor/sha_core/n3771_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3772_s7  (
	.I0(\top/processor/sha_core/n3726_139 ),
	.I1(\top/processor/sha_core/n3726_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3772_10 )
);
defparam \top/processor/sha_core/n3772_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3772_s8  (
	.I0(\top/processor/sha_core/n3726_147 ),
	.I1(\top/processor/sha_core/n3726_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3772_11 )
);
defparam \top/processor/sha_core/n3772_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3772_s9  (
	.I0(\top/processor/sha_core/n3715_139 ),
	.I1(\top/processor/sha_core/n3715_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3772_12 )
);
defparam \top/processor/sha_core/n3772_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3772_s10  (
	.I0(\top/processor/sha_core/n3715_147 ),
	.I1(\top/processor/sha_core/n3715_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3772_13 )
);
defparam \top/processor/sha_core/n3772_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3773_s7  (
	.I0(\top/processor/sha_core/n3725_139 ),
	.I1(\top/processor/sha_core/n3725_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3773_10 )
);
defparam \top/processor/sha_core/n3773_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3773_s8  (
	.I0(\top/processor/sha_core/n3725_147 ),
	.I1(\top/processor/sha_core/n3725_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3773_11 )
);
defparam \top/processor/sha_core/n3773_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3773_s9  (
	.I0(\top/processor/sha_core/n3714_139 ),
	.I1(\top/processor/sha_core/n3714_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3773_12 )
);
defparam \top/processor/sha_core/n3773_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3773_s10  (
	.I0(\top/processor/sha_core/n3714_147 ),
	.I1(\top/processor/sha_core/n3714_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3773_13 )
);
defparam \top/processor/sha_core/n3773_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3774_s7  (
	.I0(\top/processor/sha_core/n3724_139 ),
	.I1(\top/processor/sha_core/n3724_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3774_10 )
);
defparam \top/processor/sha_core/n3774_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3774_s8  (
	.I0(\top/processor/sha_core/n3724_147 ),
	.I1(\top/processor/sha_core/n3724_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3774_11 )
);
defparam \top/processor/sha_core/n3774_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3774_s9  (
	.I0(\top/processor/sha_core/n3713_139 ),
	.I1(\top/processor/sha_core/n3713_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3774_12 )
);
defparam \top/processor/sha_core/n3774_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3774_s10  (
	.I0(\top/processor/sha_core/n3713_147 ),
	.I1(\top/processor/sha_core/n3713_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3774_13 )
);
defparam \top/processor/sha_core/n3774_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3775_s7  (
	.I0(\top/processor/sha_core/n3723_135 ),
	.I1(\top/processor/sha_core/n3723_139 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3775_10 )
);
defparam \top/processor/sha_core/n3775_s7 .INIT=16'h0CFA;
LUT4 \top/processor/sha_core/n3775_s8  (
	.I0(\top/processor/sha_core/n3723_147 ),
	.I1(\top/processor/sha_core/n3723_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3775_11 )
);
defparam \top/processor/sha_core/n3775_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3775_s9  (
	.I0(\top/processor/sha_core/n3712_139 ),
	.I1(\top/processor/sha_core/n3712_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3775_12 )
);
defparam \top/processor/sha_core/n3775_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3775_s10  (
	.I0(\top/processor/sha_core/n3712_147 ),
	.I1(\top/processor/sha_core/n3712_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3775_13 )
);
defparam \top/processor/sha_core/n3775_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3776_s7  (
	.I0(\top/processor/sha_core/n3711_139 ),
	.I1(\top/processor/sha_core/n3711_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3776_10 )
);
defparam \top/processor/sha_core/n3776_s7 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3776_s8  (
	.I0(\top/processor/sha_core/n3711_147 ),
	.I1(\top/processor/sha_core/n3711_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3776_11 )
);
defparam \top/processor/sha_core/n3776_s8 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3776_s9  (
	.I0(\top/processor/sha_core/n3722_139 ),
	.I1(\top/processor/sha_core/n3722_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3776_12 )
);
defparam \top/processor/sha_core/n3776_s9 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3776_s10  (
	.I0(\top/processor/sha_core/n3722_147 ),
	.I1(\top/processor/sha_core/n3722_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3776_13 )
);
defparam \top/processor/sha_core/n3776_s10 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3777_s4  (
	.I0(\top/processor/sha_core/n3710_139 ),
	.I1(\top/processor/sha_core/n3710_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3777_7 )
);
defparam \top/processor/sha_core/n3777_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3777_s5  (
	.I0(\top/processor/sha_core/n3710_147 ),
	.I1(\top/processor/sha_core/n3710_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3777_8 )
);
defparam \top/processor/sha_core/n3777_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3778_s4  (
	.I0(\top/processor/sha_core/n3709_139 ),
	.I1(\top/processor/sha_core/n3709_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3778_7 )
);
defparam \top/processor/sha_core/n3778_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3778_s5  (
	.I0(\top/processor/sha_core/n3709_147 ),
	.I1(\top/processor/sha_core/n3709_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3778_8 )
);
defparam \top/processor/sha_core/n3778_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3779_s4  (
	.I0(\top/processor/sha_core/n3708_139 ),
	.I1(\top/processor/sha_core/n3708_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3779_7 )
);
defparam \top/processor/sha_core/n3779_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3779_s5  (
	.I0(\top/processor/sha_core/n3708_147 ),
	.I1(\top/processor/sha_core/n3708_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3779_8 )
);
defparam \top/processor/sha_core/n3779_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3780_s4  (
	.I0(\top/processor/sha_core/n3707_139 ),
	.I1(\top/processor/sha_core/n3707_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3780_7 )
);
defparam \top/processor/sha_core/n3780_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3780_s5  (
	.I0(\top/processor/sha_core/n3707_147 ),
	.I1(\top/processor/sha_core/n3707_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3780_8 )
);
defparam \top/processor/sha_core/n3780_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3781_s4  (
	.I0(\top/processor/sha_core/n3706_139 ),
	.I1(\top/processor/sha_core/n3706_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3781_7 )
);
defparam \top/processor/sha_core/n3781_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3781_s5  (
	.I0(\top/processor/sha_core/n3706_147 ),
	.I1(\top/processor/sha_core/n3706_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3781_8 )
);
defparam \top/processor/sha_core/n3781_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3782_s4  (
	.I0(\top/processor/sha_core/n3705_139 ),
	.I1(\top/processor/sha_core/n3705_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3782_7 )
);
defparam \top/processor/sha_core/n3782_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3782_s5  (
	.I0(\top/processor/sha_core/n3705_147 ),
	.I1(\top/processor/sha_core/n3705_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3782_8 )
);
defparam \top/processor/sha_core/n3782_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3783_s4  (
	.I0(\top/processor/sha_core/n3736_139 ),
	.I1(\top/processor/sha_core/n3736_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3783_7 )
);
defparam \top/processor/sha_core/n3783_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3783_s5  (
	.I0(\top/processor/sha_core/n3736_147 ),
	.I1(\top/processor/sha_core/n3736_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3783_8 )
);
defparam \top/processor/sha_core/n3783_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3784_s4  (
	.I0(\top/processor/sha_core/n3735_139 ),
	.I1(\top/processor/sha_core/n3735_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3784_7 )
);
defparam \top/processor/sha_core/n3784_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3784_s5  (
	.I0(\top/processor/sha_core/n3735_147 ),
	.I1(\top/processor/sha_core/n3735_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3784_8 )
);
defparam \top/processor/sha_core/n3784_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3785_s4  (
	.I0(\top/processor/sha_core/n3734_139 ),
	.I1(\top/processor/sha_core/n3734_135 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3785_7 )
);
defparam \top/processor/sha_core/n3785_s4 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n3785_s5  (
	.I0(\top/processor/sha_core/n3734_147 ),
	.I1(\top/processor/sha_core/n3734_143 ),
	.I2(\top/processor/sha_core/n3607_196 ),
	.I3(\top/processor/sha_core/n14441_10 ),
	.F(\top/processor/sha_core/n3785_8 )
);
defparam \top/processor/sha_core/n3785_s5 .INIT=16'hFA0C;
LUT4 \top/processor/sha_core/n8430_s11  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [95]),
	.I2(\top/processor/core_block [31]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8430_14 )
);
defparam \top/processor/sha_core/n8430_s11 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8430_s12  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [127]),
	.I2(\top/processor/core_block [63]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8430_15 )
);
defparam \top/processor/sha_core/n8430_s12 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s10  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [158]),
	.I2(\top/processor/core_block [62]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8431_13 )
);
defparam \top/processor/sha_core/n8431_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8431_s11  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [94]),
	.I2(\top/processor/core_block [30]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8431_14 )
);
defparam \top/processor/sha_core/n8431_s11 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [157]),
	.I2(\top/processor/core_block [61]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8432_12 )
);
defparam \top/processor/sha_core/n8432_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8432_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [93]),
	.I2(\top/processor/core_block [29]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8432_13 )
);
defparam \top/processor/sha_core/n8432_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [156]),
	.I2(\top/processor/core_block [60]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8433_12 )
);
defparam \top/processor/sha_core/n8433_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8433_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [92]),
	.I2(\top/processor/core_block [28]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8433_13 )
);
defparam \top/processor/sha_core/n8433_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s9  (
	.I0(\top/processor/core_block [475]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [155]),
	.I3(\top/processor/sha_core/w[11]_31_9 ),
	.F(\top/processor/sha_core/n8434_12 )
);
defparam \top/processor/sha_core/n8434_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8434_s10  (
	.I0(\top/processor/core_block [443]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [379]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8434_13 )
);
defparam \top/processor/sha_core/n8434_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s9  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [345]),
	.I2(\top/processor/core_block [89]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8436_12 )
);
defparam \top/processor/sha_core/n8436_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8436_s10  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [313]),
	.I2(\top/processor/core_block [153]),
	.I3(\top/processor/sha_core/w[11]_31_9 ),
	.F(\top/processor/sha_core/n8436_13 )
);
defparam \top/processor/sha_core/n8436_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [152]),
	.I2(\top/processor/core_block [56]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8437_12 )
);
defparam \top/processor/sha_core/n8437_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8437_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [88]),
	.I2(\top/processor/core_block [24]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8437_13 )
);
defparam \top/processor/sha_core/n8437_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s9  (
	.I0(\top/processor/core_block [503]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [279]),
	.I3(\top/processor/sha_core/w[7]_31_11 ),
	.F(\top/processor/sha_core/n8438_12 )
);
defparam \top/processor/sha_core/n8438_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8438_s10  (
	.I0(\top/processor/core_block [471]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [87]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8438_13 )
);
defparam \top/processor/sha_core/n8438_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8439_s4  (
	.I0(\top/processor/core_block [470]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [374]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8439_7 )
);
defparam \top/processor/sha_core/n8439_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8439_s5  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [502]),
	.I2(\top/processor/core_block [438]),
	.I3(\top/processor/sha_core/w[2]_31_9 ),
	.F(\top/processor/sha_core/n8439_8 )
);
defparam \top/processor/sha_core/n8439_s5 .INIT=16'h0777;
LUT3 \top/processor/sha_core/n8439_s6  (
	.I0(\top/processor/sha_core/w[15]_31_11 ),
	.I1(\top/processor/core_block [22]),
	.I2(\top/processor/sha_core/n8439_13 ),
	.F(\top/processor/sha_core/n8439_9 )
);
defparam \top/processor/sha_core/n8439_s6 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8439_s7  (
	.I0(\top/processor/sha_core/w[10]_31_9 ),
	.I1(\top/processor/core_block [182]),
	.I2(\top/processor/core_block [86]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8439_10 )
);
defparam \top/processor/sha_core/n8439_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8439_s8  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [342]),
	.I2(\top/processor/core_block [246]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8439_11 )
);
defparam \top/processor/sha_core/n8439_s8 .INIT=16'h0777;
LUT3 \top/processor/sha_core/n8439_s9  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [214]),
	.I2(\top/processor/sha_core/n8439_14 ),
	.F(\top/processor/sha_core/n8439_12 )
);
defparam \top/processor/sha_core/n8439_s9 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8440_s9  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [213]),
	.I2(\top/processor/core_block [85]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8440_12 )
);
defparam \top/processor/sha_core/n8440_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8440_s10  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [277]),
	.I2(\top/processor/core_block [245]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8440_13 )
);
defparam \top/processor/sha_core/n8440_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [148]),
	.I2(\top/processor/core_block [52]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8441_12 )
);
defparam \top/processor/sha_core/n8441_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8441_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [84]),
	.I2(\top/processor/core_block [20]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8441_13 )
);
defparam \top/processor/sha_core/n8441_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8442_s6  (
	.I0(\top/processor/core_block [371]),
	.I1(\top/processor/sha_core/w[4]_31_9 ),
	.I2(\top/processor/core_block [19]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8442_9 )
);
defparam \top/processor/sha_core/n8442_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8442_s7  (
	.I0(\top/processor/sha_core/w[6]_31_9 ),
	.I1(\top/processor/core_block [307]),
	.I2(\top/processor/core_block [179]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8442_10 )
);
defparam \top/processor/sha_core/n8442_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8442_s8  (
	.I0(\top/processor/core_block [403]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [339]),
	.I3(\top/processor/sha_core/w[5]_31_9 ),
	.F(\top/processor/sha_core/n8442_11 )
);
defparam \top/processor/sha_core/n8442_s8 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8442_s9  (
	.I0(\top/processor/core_block [499]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [275]),
	.I3(\top/processor/sha_core/w[7]_31_11 ),
	.F(\top/processor/sha_core/n8442_12 )
);
defparam \top/processor/sha_core/n8442_s9 .INIT=16'h0777;
LUT3 \top/processor/sha_core/n8442_s10  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [115]),
	.I2(\top/processor/sha_core/n8442_14 ),
	.F(\top/processor/sha_core/n8442_13 )
);
defparam \top/processor/sha_core/n8442_s10 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8443_s9  (
	.I0(\top/processor/core_block [434]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [146]),
	.I3(\top/processor/sha_core/w[11]_31_9 ),
	.F(\top/processor/sha_core/n8443_12 )
);
defparam \top/processor/sha_core/n8443_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8443_s10  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [114]),
	.I2(\top/processor/core_block [50]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8443_13 )
);
defparam \top/processor/sha_core/n8443_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s9  (
	.I0(\top/processor/core_block [465]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [337]),
	.I3(\top/processor/sha_core/w[5]_31_9 ),
	.F(\top/processor/sha_core/n8444_12 )
);
defparam \top/processor/sha_core/n8444_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8444_s10  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [497]),
	.I2(\top/processor/core_block [401]),
	.I3(\top/processor/sha_core/w[3]_31_9 ),
	.F(\top/processor/sha_core/n8444_13 )
);
defparam \top/processor/sha_core/n8444_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s9  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [79]),
	.I2(\top/processor/core_block [47]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8446_12 )
);
defparam \top/processor/sha_core/n8446_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8446_s10  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [143]),
	.I2(\top/processor/core_block [111]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8446_13 )
);
defparam \top/processor/sha_core/n8446_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s9  (
	.I0(\top/processor/core_block [398]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [142]),
	.I3(\top/processor/sha_core/w[11]_31_9 ),
	.F(\top/processor/sha_core/n8447_12 )
);
defparam \top/processor/sha_core/n8447_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8447_s10  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [334]),
	.I2(\top/processor/core_block [238]),
	.I3(\top/processor/sha_core/w[8]_31_9 ),
	.F(\top/processor/sha_core/n8447_13 )
);
defparam \top/processor/sha_core/n8447_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s9  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [205]),
	.I2(\top/processor/core_block [109]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8448_12 )
);
defparam \top/processor/sha_core/n8448_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8448_s10  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [141]),
	.I2(\top/processor/core_block [45]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8448_13 )
);
defparam \top/processor/sha_core/n8448_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s9  (
	.I0(\top/processor/core_block [492]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [172]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8449_12 )
);
defparam \top/processor/sha_core/n8449_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8449_s10  (
	.I0(\top/processor/core_block [460]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [76]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8449_13 )
);
defparam \top/processor/sha_core/n8449_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8450_s6  (
	.I0(\top/processor/core_block [427]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [363]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8450_9 )
);
defparam \top/processor/sha_core/n8450_s6 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8450_s7  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [75]),
	.I2(\top/processor/core_block [11]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8450_10 )
);
defparam \top/processor/sha_core/n8450_s7 .INIT=16'h0777;
LUT3 \top/processor/sha_core/n8450_s8  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [107]),
	.I2(\top/processor/sha_core/n8450_14 ),
	.F(\top/processor/sha_core/n8450_11 )
);
defparam \top/processor/sha_core/n8450_s8 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8450_s9  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [331]),
	.I2(\top/processor/core_block [299]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8450_12 )
);
defparam \top/processor/sha_core/n8450_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8450_s10  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [491]),
	.I2(\top/processor/core_block [459]),
	.I3(\top/processor/sha_core/n8431_6 ),
	.F(\top/processor/sha_core/n8450_13 )
);
defparam \top/processor/sha_core/n8450_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [137]),
	.I2(\top/processor/core_block [41]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8452_12 )
);
defparam \top/processor/sha_core/n8452_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8452_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [73]),
	.I2(\top/processor/core_block [9]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8452_13 )
);
defparam \top/processor/sha_core/n8452_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [136]),
	.I2(\top/processor/core_block [40]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8453_12 )
);
defparam \top/processor/sha_core/n8453_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8453_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [72]),
	.I2(\top/processor/core_block [8]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8453_13 )
);
defparam \top/processor/sha_core/n8453_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s9  (
	.I0(\top/processor/core_block [487]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [263]),
	.I3(\top/processor/sha_core/w[7]_31_11 ),
	.F(\top/processor/sha_core/n8454_12 )
);
defparam \top/processor/sha_core/n8454_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8454_s10  (
	.I0(\top/processor/core_block [455]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [71]),
	.I3(\top/processor/sha_core/w[13]_31_9 ),
	.F(\top/processor/sha_core/n8454_13 )
);
defparam \top/processor/sha_core/n8454_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s9  (
	.I0(\top/processor/core_block [421]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [389]),
	.I3(\top/processor/sha_core/w[3]_31_9 ),
	.F(\top/processor/sha_core/n8456_12 )
);
defparam \top/processor/sha_core/n8456_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8456_s10  (
	.I0(\top/processor/core_block [485]),
	.I1(\top/processor/sha_core/n8430_11 ),
	.I2(\top/processor/core_block [357]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8456_13 )
);
defparam \top/processor/sha_core/n8456_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8457_s4  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [260]),
	.I2(\top/processor/core_block [164]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8457_7 )
);
defparam \top/processor/sha_core/n8457_s4 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8457_s5  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [68]),
	.I2(\top/processor/core_block [4]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8457_8 )
);
defparam \top/processor/sha_core/n8457_s5 .INIT=16'h0777;
LUT3 \top/processor/sha_core/n8457_s6  (
	.I0(\top/processor/sha_core/w[3]_31_9 ),
	.I1(\top/processor/core_block [388]),
	.I2(\top/processor/sha_core/n8457_12 ),
	.F(\top/processor/sha_core/n8457_9 )
);
defparam \top/processor/sha_core/n8457_s6 .INIT=8'h70;
LUT4 \top/processor/sha_core/n8457_s7  (
	.I0(\top/processor/sha_core/w[5]_31_9 ),
	.I1(\top/processor/core_block [324]),
	.I2(\top/processor/core_block [292]),
	.I3(\top/processor/sha_core/w[6]_31_9 ),
	.F(\top/processor/sha_core/n8457_10 )
);
defparam \top/processor/sha_core/n8457_s7 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8457_s8  (
	.I0(\top/processor/sha_core/n8430_11 ),
	.I1(\top/processor/core_block [484]),
	.I2(\top/processor/sha_core/n8457_13 ),
	.I3(\top/processor/sha_core/n8457_14 ),
	.F(\top/processor/sha_core/n8457_11 )
);
defparam \top/processor/sha_core/n8457_s8 .INIT=16'h7000;
LUT4 \top/processor/sha_core/n8458_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [131]),
	.I2(\top/processor/core_block [35]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8458_12 )
);
defparam \top/processor/sha_core/n8458_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8458_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [67]),
	.I2(\top/processor/core_block [3]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8458_13 )
);
defparam \top/processor/sha_core/n8458_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s9  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [130]),
	.I2(\top/processor/core_block [34]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8459_12 )
);
defparam \top/processor/sha_core/n8459_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8459_s10  (
	.I0(\top/processor/sha_core/w[13]_31_9 ),
	.I1(\top/processor/core_block [66]),
	.I2(\top/processor/core_block [2]),
	.I3(\top/processor/sha_core/w[15]_31_11 ),
	.F(\top/processor/sha_core/n8459_13 )
);
defparam \top/processor/sha_core/n8459_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s9  (
	.I0(\top/processor/core_block [385]),
	.I1(\top/processor/sha_core/w[3]_31_9 ),
	.I2(\top/processor/core_block [193]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8460_12 )
);
defparam \top/processor/sha_core/n8460_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8460_s10  (
	.I0(\top/processor/core_block [417]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [97]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8460_13 )
);
defparam \top/processor/sha_core/n8460_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s9  (
	.I0(\top/processor/sha_core/w[9]_31_9 ),
	.I1(\top/processor/core_block [192]),
	.I2(\top/processor/core_block [96]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8461_12 )
);
defparam \top/processor/sha_core/n8461_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8461_s10  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [256]),
	.I2(\top/processor/core_block [160]),
	.I3(\top/processor/sha_core/w[10]_31_9 ),
	.F(\top/processor/sha_core/n8461_13 )
);
defparam \top/processor/sha_core/n8461_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8439_s10  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [150]),
	.I2(\top/processor/core_block [54]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8439_13 )
);
defparam \top/processor/sha_core/n8439_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8439_s11  (
	.I0(\top/processor/sha_core/w[7]_31_11 ),
	.I1(\top/processor/core_block [278]),
	.I2(\top/processor/core_block [118]),
	.I3(\top/processor/sha_core/w[12]_31_9 ),
	.F(\top/processor/sha_core/n8439_14 )
);
defparam \top/processor/sha_core/n8439_s11 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8442_s11  (
	.I0(\top/processor/core_block [435]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [211]),
	.I3(\top/processor/sha_core/w[9]_31_9 ),
	.F(\top/processor/sha_core/n8442_14 )
);
defparam \top/processor/sha_core/n8442_s11 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8450_s11  (
	.I0(\top/processor/sha_core/w[11]_31_9 ),
	.I1(\top/processor/core_block [139]),
	.I2(\top/processor/core_block [43]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8450_14 )
);
defparam \top/processor/sha_core/n8450_s11 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8457_s9  (
	.I0(\top/processor/core_block [452]),
	.I1(\top/processor/sha_core/n8431_6 ),
	.I2(\top/processor/core_block [356]),
	.I3(\top/processor/sha_core/w[4]_31_9 ),
	.F(\top/processor/sha_core/n8457_12 )
);
defparam \top/processor/sha_core/n8457_s9 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8457_s10  (
	.I0(\top/processor/core_block [420]),
	.I1(\top/processor/sha_core/w[2]_31_9 ),
	.I2(\top/processor/core_block [132]),
	.I3(\top/processor/sha_core/w[11]_31_9 ),
	.F(\top/processor/sha_core/n8457_13 )
);
defparam \top/processor/sha_core/n8457_s10 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n8457_s11  (
	.I0(\top/processor/sha_core/w[12]_31_9 ),
	.I1(\top/processor/core_block [100]),
	.I2(\top/processor/core_block [36]),
	.I3(\top/processor/sha_core/w[14]_31_9 ),
	.F(\top/processor/sha_core/n8457_14 )
);
defparam \top/processor/sha_core/n8457_s11 .INIT=16'h0777;
LUT4 \top/processor/sha_core/n293_s5813  (
	.I0(\top/processor/sha_core/t [4]),
	.I1(\top/processor/sha_core/t [5]),
	.I2(\top/processor/sha_core/t [2]),
	.I3(\top/processor/sha_core/t [3]),
	.F(\top/processor/sha_core/n293_7386 )
);
defparam \top/processor/sha_core/n293_s5813 .INIT=16'h1055;
LUT4 \top/processor/sha_core/n293_s5814  (
	.I0(\top/processor/sha_core/t [2]),
	.I1(\top/processor/sha_core/t [3]),
	.I2(\top/processor/sha_core/t [4]),
	.I3(\top/processor/sha_core/t [5]),
	.F(\top/processor/sha_core/n293_7388 )
);
defparam \top/processor/sha_core/n293_s5814 .INIT=16'hBACF;
LUT4 \top/processor/sha_core/n3766_s12  (
	.I0(\top/processor/sha_core/n3766_6 ),
	.I1(\top/processor/sha_core/n3766_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.I3(\top/processor/sha_core/n3766_5 ),
	.F(\top/processor/sha_core/n3766_16 )
);
defparam \top/processor/sha_core/n3766_s12 .INIT=16'h53AC;
LUT4 \top/processor/sha_core/n3767_s11  (
	.I0(\top/processor/sha_core/n3767_6 ),
	.I1(\top/processor/sha_core/n3767_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.I3(\top/processor/sha_core/n3767_5 ),
	.F(\top/processor/sha_core/n3767_15 )
);
defparam \top/processor/sha_core/n3767_s11 .INIT=16'h53AC;
LUT4 \top/processor/sha_core/n3768_s11  (
	.I0(\top/processor/sha_core/n3768_6 ),
	.I1(\top/processor/sha_core/n3768_7 ),
	.I2(\top/processor/sha_core/n3766_8 ),
	.I3(\top/processor/sha_core/n3768_5 ),
	.F(\top/processor/sha_core/n3768_15 )
);
defparam \top/processor/sha_core/n3768_s11 .INIT=16'h53AC;
LUT4 \top/processor/sha_core/n3607_s167  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.I3(\top/processor/sha_core/msg_idx [2]),
	.F(\top/processor/sha_core/n3607_196 )
);
defparam \top/processor/sha_core/n3607_s167 .INIT=16'h9555;
LUT4 \top/processor/sha_core/w[31]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [3]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.I3(\top/processor/sha_core/msg_idx [2]),
	.F(\top/processor/sha_core/w[31]_31_11 )
);
defparam \top/processor/sha_core/w[31]_31_s6 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[23]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[63]_31_9 ),
	.F(\top/processor/sha_core/w[23]_31_11 )
);
defparam \top/processor/sha_core/w[23]_31_s6 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[15]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[40]_31_9 ),
	.F(\top/processor/sha_core/w[15]_31_11 )
);
defparam \top/processor/sha_core/w[15]_31_s6 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[7]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [1]),
	.I1(\top/processor/sha_core/msg_idx [0]),
	.I2(\top/processor/sha_core/msg_idx [2]),
	.I3(\top/processor/sha_core/w[0]_31_9 ),
	.F(\top/processor/sha_core/w[7]_31_11 )
);
defparam \top/processor/sha_core/w[7]_31_s6 .INIT=16'h8000;
LUT4 \top/processor/sha_core/w[2]_31_s7  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [6]),
	.I2(\top/processor/sha_core/state [1]),
	.I3(\top/processor/sha_core/state [0]),
	.F(\top/processor/sha_core/w[2]_31_12 )
);
defparam \top/processor/sha_core/w[2]_31_s7 .INIT=16'h0100;
LUT4 \top/processor/sha_core/w[47]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[23]_31_11 ),
	.F(\top/processor/sha_core/w[47]_31_10 )
);
defparam \top/processor/sha_core/w[47]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[46]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[22]_31_9 ),
	.F(\top/processor/sha_core/w[46]_31_10 )
);
defparam \top/processor/sha_core/w[46]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[45]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[21]_31_9 ),
	.F(\top/processor/sha_core/w[45]_31_10 )
);
defparam \top/processor/sha_core/w[45]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[44]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[20]_31_9 ),
	.F(\top/processor/sha_core/w[44]_31_10 )
);
defparam \top/processor/sha_core/w[44]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[43]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[19]_31_9 ),
	.F(\top/processor/sha_core/w[43]_31_10 )
);
defparam \top/processor/sha_core/w[43]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[42]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[18]_31_9 ),
	.F(\top/processor/sha_core/w[42]_31_10 )
);
defparam \top/processor/sha_core/w[42]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[41]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[41]_31_10 )
);
defparam \top/processor/sha_core/w[41]_31_s5 .INIT=16'h2000;
LUT4 \top/processor/sha_core/w[40]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[40]_31_11 )
);
defparam \top/processor/sha_core/w[40]_31_s6 .INIT=16'h2000;
LUT4 \top/processor/sha_core/n3577_s4  (
	.I0(\top/processor/sha_core/n3578_12 ),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/msg_idx [5]),
	.F(\top/processor/sha_core/n3577_11 )
);
defparam \top/processor/sha_core/n3577_s4 .INIT=16'hFE01;
LUT4 \top/processor/sha_core/w[39]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[23]_31_11 ),
	.F(\top/processor/sha_core/w[39]_31_10 )
);
defparam \top/processor/sha_core/w[39]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[38]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[22]_31_9 ),
	.F(\top/processor/sha_core/w[38]_31_10 )
);
defparam \top/processor/sha_core/w[38]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[37]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[21]_31_9 ),
	.F(\top/processor/sha_core/w[37]_31_10 )
);
defparam \top/processor/sha_core/w[37]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[36]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[20]_31_9 ),
	.F(\top/processor/sha_core/w[36]_31_10 )
);
defparam \top/processor/sha_core/w[36]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[35]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[19]_31_9 ),
	.F(\top/processor/sha_core/w[35]_31_10 )
);
defparam \top/processor/sha_core/w[35]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[34]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[18]_31_9 ),
	.F(\top/processor/sha_core/w[34]_31_10 )
);
defparam \top/processor/sha_core/w[34]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[33]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[33]_31_10 )
);
defparam \top/processor/sha_core/w[33]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[32]_31_s5  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[32]_31_10 )
);
defparam \top/processor/sha_core/w[32]_31_s5 .INIT=16'h0200;
LUT4 \top/processor/sha_core/w[1]_31_s6  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[1]_31_9 ),
	.F(\top/processor/sha_core/w[1]_31_11 )
);
defparam \top/processor/sha_core/w[1]_31_s6 .INIT=16'h0100;
LUT4 \top/processor/sha_core/w[0]_31_s7  (
	.I0(\top/processor/sha_core/msg_idx [5]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/msg_idx [3]),
	.I3(\top/processor/sha_core/w[0]_31_10 ),
	.F(\top/processor/sha_core/w[0]_31_12 )
);
defparam \top/processor/sha_core/w[0]_31_s7 .INIT=16'h0100;
LUT3 \top/processor/sha_core/n14441_s6  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/msg_idx [4]),
	.I2(\top/processor/sha_core/w[31]_31_11 ),
	.F(\top/processor/sha_core/n14441_12 )
);
defparam \top/processor/sha_core/n14441_s6 .INIT=8'h28;
LUT4 \top/processor/sha_core/n14443_s5  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.I3(\top/processor/sha_core/msg_idx [2]),
	.F(\top/processor/sha_core/n14443_11 )
);
defparam \top/processor/sha_core/n14443_s5 .INIT=16'h2A80;
LUT3 \top/processor/sha_core/n14444_s5  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/msg_idx [1]),
	.I2(\top/processor/sha_core/msg_idx [0]),
	.F(\top/processor/sha_core/n14444_11 )
);
defparam \top/processor/sha_core/n14444_s5 .INIT=8'h28;
LUT4 \top/processor/sha_core/n3544_s1  (
	.I0(\top/processor/sha_core/n3510_189 ),
	.I1(\top/processor/sha_core/n3510_191 ),
	.I2(\top/processor/sha_core/n3459_9 ),
	.I3(\top/processor/sha_core/n3508_193 ),
	.F(\top/processor/sha_core/n3544_5 )
);
defparam \top/processor/sha_core/n3544_s1 .INIT=16'h35CA;
LUT4 \top/processor/sha_core/n3542_s1  (
	.I0(\top/processor/sha_core/n3512_193 ),
	.I1(\top/processor/sha_core/n3510_189 ),
	.I2(\top/processor/sha_core/n3510_191 ),
	.I3(\top/processor/sha_core/n3459_9 ),
	.F(\top/processor/sha_core/n3542_5 )
);
defparam \top/processor/sha_core/n3542_s1 .INIT=16'h5A66;
LUT4 \top/processor/sha_core/n11871_s8  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/state_0_9 ),
	.I2(\top/processor/core_start ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11871_15 )
);
defparam \top/processor/sha_core/n11871_s8 .INIT=16'hE4D8;
LUT4 \top/processor/sha_core/n11870_s8  (
	.I0(\top/processor/sha_core/state [0]),
	.I1(\top/processor/sha_core/state_0_9 ),
	.I2(\top/processor/core_start ),
	.I3(\top/processor/sha_core/state [1]),
	.F(\top/processor/sha_core/n11870_15 )
);
defparam \top/processor/sha_core/n11870_s8 .INIT=16'hF522;
DFFCE \top/processor/sha_core/hash_out_255_s0  (
	.D(\top/processor/sha_core/h0 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [255])
);
defparam \top/processor/sha_core/hash_out_255_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_254_s0  (
	.D(\top/processor/sha_core/h0 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [254])
);
defparam \top/processor/sha_core/hash_out_254_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_253_s0  (
	.D(\top/processor/sha_core/h0 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [253])
);
defparam \top/processor/sha_core/hash_out_253_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_252_s0  (
	.D(\top/processor/sha_core/h0 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [252])
);
defparam \top/processor/sha_core/hash_out_252_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_251_s0  (
	.D(\top/processor/sha_core/h0 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [251])
);
defparam \top/processor/sha_core/hash_out_251_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_250_s0  (
	.D(\top/processor/sha_core/h0 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [250])
);
defparam \top/processor/sha_core/hash_out_250_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_249_s0  (
	.D(\top/processor/sha_core/h0 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [249])
);
defparam \top/processor/sha_core/hash_out_249_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_248_s0  (
	.D(\top/processor/sha_core/h0 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [248])
);
defparam \top/processor/sha_core/hash_out_248_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_247_s0  (
	.D(\top/processor/sha_core/h0 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [247])
);
defparam \top/processor/sha_core/hash_out_247_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_246_s0  (
	.D(\top/processor/sha_core/h0 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [246])
);
defparam \top/processor/sha_core/hash_out_246_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_245_s0  (
	.D(\top/processor/sha_core/h0 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [245])
);
defparam \top/processor/sha_core/hash_out_245_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_244_s0  (
	.D(\top/processor/sha_core/h0 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [244])
);
defparam \top/processor/sha_core/hash_out_244_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_243_s0  (
	.D(\top/processor/sha_core/h0 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [243])
);
defparam \top/processor/sha_core/hash_out_243_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_242_s0  (
	.D(\top/processor/sha_core/h0 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [242])
);
defparam \top/processor/sha_core/hash_out_242_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_241_s0  (
	.D(\top/processor/sha_core/h0 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [241])
);
defparam \top/processor/sha_core/hash_out_241_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_240_s0  (
	.D(\top/processor/sha_core/h0 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [240])
);
defparam \top/processor/sha_core/hash_out_240_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_239_s0  (
	.D(\top/processor/sha_core/h0 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [239])
);
defparam \top/processor/sha_core/hash_out_239_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_238_s0  (
	.D(\top/processor/sha_core/h0 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [238])
);
defparam \top/processor/sha_core/hash_out_238_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_237_s0  (
	.D(\top/processor/sha_core/h0 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [237])
);
defparam \top/processor/sha_core/hash_out_237_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_236_s0  (
	.D(\top/processor/sha_core/h0 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [236])
);
defparam \top/processor/sha_core/hash_out_236_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_235_s0  (
	.D(\top/processor/sha_core/h0 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [235])
);
defparam \top/processor/sha_core/hash_out_235_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_234_s0  (
	.D(\top/processor/sha_core/h0 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [234])
);
defparam \top/processor/sha_core/hash_out_234_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_233_s0  (
	.D(\top/processor/sha_core/h0 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [233])
);
defparam \top/processor/sha_core/hash_out_233_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_232_s0  (
	.D(\top/processor/sha_core/h0 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [232])
);
defparam \top/processor/sha_core/hash_out_232_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_231_s0  (
	.D(\top/processor/sha_core/h0 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [231])
);
defparam \top/processor/sha_core/hash_out_231_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_230_s0  (
	.D(\top/processor/sha_core/h0 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [230])
);
defparam \top/processor/sha_core/hash_out_230_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_229_s0  (
	.D(\top/processor/sha_core/h0 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [229])
);
defparam \top/processor/sha_core/hash_out_229_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_228_s0  (
	.D(\top/processor/sha_core/h0 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [228])
);
defparam \top/processor/sha_core/hash_out_228_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_227_s0  (
	.D(\top/processor/sha_core/h0 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [227])
);
defparam \top/processor/sha_core/hash_out_227_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_226_s0  (
	.D(\top/processor/sha_core/h0 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [226])
);
defparam \top/processor/sha_core/hash_out_226_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_225_s0  (
	.D(\top/processor/sha_core/h0 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [225])
);
defparam \top/processor/sha_core/hash_out_225_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_224_s0  (
	.D(\top/processor/sha_core/h0 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [224])
);
defparam \top/processor/sha_core/hash_out_224_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_223_s0  (
	.D(\top/processor/sha_core/h1 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [223])
);
defparam \top/processor/sha_core/hash_out_223_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_222_s0  (
	.D(\top/processor/sha_core/h1 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [222])
);
defparam \top/processor/sha_core/hash_out_222_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_221_s0  (
	.D(\top/processor/sha_core/h1 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [221])
);
defparam \top/processor/sha_core/hash_out_221_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_220_s0  (
	.D(\top/processor/sha_core/h1 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [220])
);
defparam \top/processor/sha_core/hash_out_220_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_219_s0  (
	.D(\top/processor/sha_core/h1 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [219])
);
defparam \top/processor/sha_core/hash_out_219_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_218_s0  (
	.D(\top/processor/sha_core/h1 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [218])
);
defparam \top/processor/sha_core/hash_out_218_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_217_s0  (
	.D(\top/processor/sha_core/h1 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [217])
);
defparam \top/processor/sha_core/hash_out_217_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_216_s0  (
	.D(\top/processor/sha_core/h1 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [216])
);
defparam \top/processor/sha_core/hash_out_216_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_215_s0  (
	.D(\top/processor/sha_core/h1 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [215])
);
defparam \top/processor/sha_core/hash_out_215_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_214_s0  (
	.D(\top/processor/sha_core/h1 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [214])
);
defparam \top/processor/sha_core/hash_out_214_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_213_s0  (
	.D(\top/processor/sha_core/h1 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [213])
);
defparam \top/processor/sha_core/hash_out_213_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_212_s0  (
	.D(\top/processor/sha_core/h1 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [212])
);
defparam \top/processor/sha_core/hash_out_212_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_211_s0  (
	.D(\top/processor/sha_core/h1 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [211])
);
defparam \top/processor/sha_core/hash_out_211_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_210_s0  (
	.D(\top/processor/sha_core/h1 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [210])
);
defparam \top/processor/sha_core/hash_out_210_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_209_s0  (
	.D(\top/processor/sha_core/h1 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [209])
);
defparam \top/processor/sha_core/hash_out_209_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_208_s0  (
	.D(\top/processor/sha_core/h1 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [208])
);
defparam \top/processor/sha_core/hash_out_208_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_207_s0  (
	.D(\top/processor/sha_core/h1 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [207])
);
defparam \top/processor/sha_core/hash_out_207_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_206_s0  (
	.D(\top/processor/sha_core/h1 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [206])
);
defparam \top/processor/sha_core/hash_out_206_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_205_s0  (
	.D(\top/processor/sha_core/h1 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [205])
);
defparam \top/processor/sha_core/hash_out_205_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_204_s0  (
	.D(\top/processor/sha_core/h1 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [204])
);
defparam \top/processor/sha_core/hash_out_204_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_203_s0  (
	.D(\top/processor/sha_core/h1 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [203])
);
defparam \top/processor/sha_core/hash_out_203_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_202_s0  (
	.D(\top/processor/sha_core/h1 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [202])
);
defparam \top/processor/sha_core/hash_out_202_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_201_s0  (
	.D(\top/processor/sha_core/h1 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [201])
);
defparam \top/processor/sha_core/hash_out_201_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_200_s0  (
	.D(\top/processor/sha_core/h1 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [200])
);
defparam \top/processor/sha_core/hash_out_200_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_199_s0  (
	.D(\top/processor/sha_core/h1 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [199])
);
defparam \top/processor/sha_core/hash_out_199_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_198_s0  (
	.D(\top/processor/sha_core/h1 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [198])
);
defparam \top/processor/sha_core/hash_out_198_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_197_s0  (
	.D(\top/processor/sha_core/h1 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [197])
);
defparam \top/processor/sha_core/hash_out_197_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_196_s0  (
	.D(\top/processor/sha_core/h1 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [196])
);
defparam \top/processor/sha_core/hash_out_196_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_195_s0  (
	.D(\top/processor/sha_core/h1 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [195])
);
defparam \top/processor/sha_core/hash_out_195_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_194_s0  (
	.D(\top/processor/sha_core/h1 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [194])
);
defparam \top/processor/sha_core/hash_out_194_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_193_s0  (
	.D(\top/processor/sha_core/h1 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [193])
);
defparam \top/processor/sha_core/hash_out_193_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_192_s0  (
	.D(\top/processor/sha_core/h1 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [192])
);
defparam \top/processor/sha_core/hash_out_192_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_191_s0  (
	.D(\top/processor/sha_core/h2 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [191])
);
defparam \top/processor/sha_core/hash_out_191_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_190_s0  (
	.D(\top/processor/sha_core/h2 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [190])
);
defparam \top/processor/sha_core/hash_out_190_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_189_s0  (
	.D(\top/processor/sha_core/h2 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [189])
);
defparam \top/processor/sha_core/hash_out_189_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_188_s0  (
	.D(\top/processor/sha_core/h2 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [188])
);
defparam \top/processor/sha_core/hash_out_188_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_187_s0  (
	.D(\top/processor/sha_core/h2 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [187])
);
defparam \top/processor/sha_core/hash_out_187_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_186_s0  (
	.D(\top/processor/sha_core/h2 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [186])
);
defparam \top/processor/sha_core/hash_out_186_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_185_s0  (
	.D(\top/processor/sha_core/h2 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [185])
);
defparam \top/processor/sha_core/hash_out_185_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_184_s0  (
	.D(\top/processor/sha_core/h2 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [184])
);
defparam \top/processor/sha_core/hash_out_184_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_183_s0  (
	.D(\top/processor/sha_core/h2 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [183])
);
defparam \top/processor/sha_core/hash_out_183_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_182_s0  (
	.D(\top/processor/sha_core/h2 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [182])
);
defparam \top/processor/sha_core/hash_out_182_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_181_s0  (
	.D(\top/processor/sha_core/h2 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [181])
);
defparam \top/processor/sha_core/hash_out_181_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_180_s0  (
	.D(\top/processor/sha_core/h2 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [180])
);
defparam \top/processor/sha_core/hash_out_180_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_179_s0  (
	.D(\top/processor/sha_core/h2 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [179])
);
defparam \top/processor/sha_core/hash_out_179_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_178_s0  (
	.D(\top/processor/sha_core/h2 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [178])
);
defparam \top/processor/sha_core/hash_out_178_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_177_s0  (
	.D(\top/processor/sha_core/h2 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [177])
);
defparam \top/processor/sha_core/hash_out_177_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_176_s0  (
	.D(\top/processor/sha_core/h2 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [176])
);
defparam \top/processor/sha_core/hash_out_176_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_175_s0  (
	.D(\top/processor/sha_core/h2 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [175])
);
defparam \top/processor/sha_core/hash_out_175_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_174_s0  (
	.D(\top/processor/sha_core/h2 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [174])
);
defparam \top/processor/sha_core/hash_out_174_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_173_s0  (
	.D(\top/processor/sha_core/h2 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [173])
);
defparam \top/processor/sha_core/hash_out_173_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_172_s0  (
	.D(\top/processor/sha_core/h2 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [172])
);
defparam \top/processor/sha_core/hash_out_172_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_171_s0  (
	.D(\top/processor/sha_core/h2 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [171])
);
defparam \top/processor/sha_core/hash_out_171_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_170_s0  (
	.D(\top/processor/sha_core/h2 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [170])
);
defparam \top/processor/sha_core/hash_out_170_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_169_s0  (
	.D(\top/processor/sha_core/h2 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [169])
);
defparam \top/processor/sha_core/hash_out_169_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_168_s0  (
	.D(\top/processor/sha_core/h2 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [168])
);
defparam \top/processor/sha_core/hash_out_168_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_167_s0  (
	.D(\top/processor/sha_core/h2 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [167])
);
defparam \top/processor/sha_core/hash_out_167_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_166_s0  (
	.D(\top/processor/sha_core/h2 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [166])
);
defparam \top/processor/sha_core/hash_out_166_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_165_s0  (
	.D(\top/processor/sha_core/h2 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [165])
);
defparam \top/processor/sha_core/hash_out_165_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_164_s0  (
	.D(\top/processor/sha_core/h2 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [164])
);
defparam \top/processor/sha_core/hash_out_164_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_163_s0  (
	.D(\top/processor/sha_core/h2 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [163])
);
defparam \top/processor/sha_core/hash_out_163_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_162_s0  (
	.D(\top/processor/sha_core/h2 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [162])
);
defparam \top/processor/sha_core/hash_out_162_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_161_s0  (
	.D(\top/processor/sha_core/h2 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [161])
);
defparam \top/processor/sha_core/hash_out_161_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_160_s0  (
	.D(\top/processor/sha_core/h2 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [160])
);
defparam \top/processor/sha_core/hash_out_160_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_159_s0  (
	.D(\top/processor/sha_core/h3 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [159])
);
defparam \top/processor/sha_core/hash_out_159_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_158_s0  (
	.D(\top/processor/sha_core/h3 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [158])
);
defparam \top/processor/sha_core/hash_out_158_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_157_s0  (
	.D(\top/processor/sha_core/h3 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [157])
);
defparam \top/processor/sha_core/hash_out_157_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_156_s0  (
	.D(\top/processor/sha_core/h3 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [156])
);
defparam \top/processor/sha_core/hash_out_156_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_155_s0  (
	.D(\top/processor/sha_core/h3 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [155])
);
defparam \top/processor/sha_core/hash_out_155_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_154_s0  (
	.D(\top/processor/sha_core/h3 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [154])
);
defparam \top/processor/sha_core/hash_out_154_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_153_s0  (
	.D(\top/processor/sha_core/h3 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [153])
);
defparam \top/processor/sha_core/hash_out_153_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_152_s0  (
	.D(\top/processor/sha_core/h3 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [152])
);
defparam \top/processor/sha_core/hash_out_152_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_151_s0  (
	.D(\top/processor/sha_core/h3 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [151])
);
defparam \top/processor/sha_core/hash_out_151_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_150_s0  (
	.D(\top/processor/sha_core/h3 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [150])
);
defparam \top/processor/sha_core/hash_out_150_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_149_s0  (
	.D(\top/processor/sha_core/h3 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [149])
);
defparam \top/processor/sha_core/hash_out_149_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_148_s0  (
	.D(\top/processor/sha_core/h3 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [148])
);
defparam \top/processor/sha_core/hash_out_148_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_147_s0  (
	.D(\top/processor/sha_core/h3 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [147])
);
defparam \top/processor/sha_core/hash_out_147_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_146_s0  (
	.D(\top/processor/sha_core/h3 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [146])
);
defparam \top/processor/sha_core/hash_out_146_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_145_s0  (
	.D(\top/processor/sha_core/h3 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [145])
);
defparam \top/processor/sha_core/hash_out_145_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_144_s0  (
	.D(\top/processor/sha_core/h3 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [144])
);
defparam \top/processor/sha_core/hash_out_144_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_143_s0  (
	.D(\top/processor/sha_core/h3 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [143])
);
defparam \top/processor/sha_core/hash_out_143_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_142_s0  (
	.D(\top/processor/sha_core/h3 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [142])
);
defparam \top/processor/sha_core/hash_out_142_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_141_s0  (
	.D(\top/processor/sha_core/h3 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [141])
);
defparam \top/processor/sha_core/hash_out_141_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_140_s0  (
	.D(\top/processor/sha_core/h3 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [140])
);
defparam \top/processor/sha_core/hash_out_140_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_139_s0  (
	.D(\top/processor/sha_core/h3 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [139])
);
defparam \top/processor/sha_core/hash_out_139_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_138_s0  (
	.D(\top/processor/sha_core/h3 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [138])
);
defparam \top/processor/sha_core/hash_out_138_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_137_s0  (
	.D(\top/processor/sha_core/h3 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [137])
);
defparam \top/processor/sha_core/hash_out_137_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_136_s0  (
	.D(\top/processor/sha_core/h3 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [136])
);
defparam \top/processor/sha_core/hash_out_136_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_135_s0  (
	.D(\top/processor/sha_core/h3 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [135])
);
defparam \top/processor/sha_core/hash_out_135_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_134_s0  (
	.D(\top/processor/sha_core/h3 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [134])
);
defparam \top/processor/sha_core/hash_out_134_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_133_s0  (
	.D(\top/processor/sha_core/h3 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [133])
);
defparam \top/processor/sha_core/hash_out_133_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_132_s0  (
	.D(\top/processor/sha_core/h3 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [132])
);
defparam \top/processor/sha_core/hash_out_132_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_131_s0  (
	.D(\top/processor/sha_core/h3 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [131])
);
defparam \top/processor/sha_core/hash_out_131_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_130_s0  (
	.D(\top/processor/sha_core/h3 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [130])
);
defparam \top/processor/sha_core/hash_out_130_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_129_s0  (
	.D(\top/processor/sha_core/h3 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [129])
);
defparam \top/processor/sha_core/hash_out_129_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_128_s0  (
	.D(\top/processor/sha_core/h3 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [128])
);
defparam \top/processor/sha_core/hash_out_128_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_127_s0  (
	.D(\top/processor/sha_core/h4 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [127])
);
defparam \top/processor/sha_core/hash_out_127_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_126_s0  (
	.D(\top/processor/sha_core/h4 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [126])
);
defparam \top/processor/sha_core/hash_out_126_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_125_s0  (
	.D(\top/processor/sha_core/h4 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [125])
);
defparam \top/processor/sha_core/hash_out_125_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_124_s0  (
	.D(\top/processor/sha_core/h4 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [124])
);
defparam \top/processor/sha_core/hash_out_124_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_123_s0  (
	.D(\top/processor/sha_core/h4 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [123])
);
defparam \top/processor/sha_core/hash_out_123_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_122_s0  (
	.D(\top/processor/sha_core/h4 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [122])
);
defparam \top/processor/sha_core/hash_out_122_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_121_s0  (
	.D(\top/processor/sha_core/h4 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [121])
);
defparam \top/processor/sha_core/hash_out_121_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_120_s0  (
	.D(\top/processor/sha_core/h4 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [120])
);
defparam \top/processor/sha_core/hash_out_120_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_119_s0  (
	.D(\top/processor/sha_core/h4 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [119])
);
defparam \top/processor/sha_core/hash_out_119_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_118_s0  (
	.D(\top/processor/sha_core/h4 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [118])
);
defparam \top/processor/sha_core/hash_out_118_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_117_s0  (
	.D(\top/processor/sha_core/h4 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [117])
);
defparam \top/processor/sha_core/hash_out_117_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_116_s0  (
	.D(\top/processor/sha_core/h4 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [116])
);
defparam \top/processor/sha_core/hash_out_116_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_115_s0  (
	.D(\top/processor/sha_core/h4 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [115])
);
defparam \top/processor/sha_core/hash_out_115_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_114_s0  (
	.D(\top/processor/sha_core/h4 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [114])
);
defparam \top/processor/sha_core/hash_out_114_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_113_s0  (
	.D(\top/processor/sha_core/h4 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [113])
);
defparam \top/processor/sha_core/hash_out_113_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_112_s0  (
	.D(\top/processor/sha_core/h4 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [112])
);
defparam \top/processor/sha_core/hash_out_112_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_111_s0  (
	.D(\top/processor/sha_core/h4 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [111])
);
defparam \top/processor/sha_core/hash_out_111_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_110_s0  (
	.D(\top/processor/sha_core/h4 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [110])
);
defparam \top/processor/sha_core/hash_out_110_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_109_s0  (
	.D(\top/processor/sha_core/h4 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [109])
);
defparam \top/processor/sha_core/hash_out_109_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_108_s0  (
	.D(\top/processor/sha_core/h4 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [108])
);
defparam \top/processor/sha_core/hash_out_108_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_107_s0  (
	.D(\top/processor/sha_core/h4 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [107])
);
defparam \top/processor/sha_core/hash_out_107_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_106_s0  (
	.D(\top/processor/sha_core/h4 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [106])
);
defparam \top/processor/sha_core/hash_out_106_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_105_s0  (
	.D(\top/processor/sha_core/h4 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [105])
);
defparam \top/processor/sha_core/hash_out_105_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_104_s0  (
	.D(\top/processor/sha_core/h4 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [104])
);
defparam \top/processor/sha_core/hash_out_104_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_103_s0  (
	.D(\top/processor/sha_core/h4 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [103])
);
defparam \top/processor/sha_core/hash_out_103_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_102_s0  (
	.D(\top/processor/sha_core/h4 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [102])
);
defparam \top/processor/sha_core/hash_out_102_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_101_s0  (
	.D(\top/processor/sha_core/h4 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [101])
);
defparam \top/processor/sha_core/hash_out_101_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_100_s0  (
	.D(\top/processor/sha_core/h4 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [100])
);
defparam \top/processor/sha_core/hash_out_100_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_99_s0  (
	.D(\top/processor/sha_core/h4 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [99])
);
defparam \top/processor/sha_core/hash_out_99_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_98_s0  (
	.D(\top/processor/sha_core/h4 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [98])
);
defparam \top/processor/sha_core/hash_out_98_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_97_s0  (
	.D(\top/processor/sha_core/h4 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [97])
);
defparam \top/processor/sha_core/hash_out_97_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_96_s0  (
	.D(\top/processor/sha_core/h4 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [96])
);
defparam \top/processor/sha_core/hash_out_96_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_95_s0  (
	.D(\top/processor/sha_core/h5 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [95])
);
defparam \top/processor/sha_core/hash_out_95_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_94_s0  (
	.D(\top/processor/sha_core/h5 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [94])
);
defparam \top/processor/sha_core/hash_out_94_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_93_s0  (
	.D(\top/processor/sha_core/h5 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [93])
);
defparam \top/processor/sha_core/hash_out_93_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_92_s0  (
	.D(\top/processor/sha_core/h5 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [92])
);
defparam \top/processor/sha_core/hash_out_92_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_91_s0  (
	.D(\top/processor/sha_core/h5 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [91])
);
defparam \top/processor/sha_core/hash_out_91_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_90_s0  (
	.D(\top/processor/sha_core/h5 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [90])
);
defparam \top/processor/sha_core/hash_out_90_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_89_s0  (
	.D(\top/processor/sha_core/h5 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [89])
);
defparam \top/processor/sha_core/hash_out_89_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_88_s0  (
	.D(\top/processor/sha_core/h5 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [88])
);
defparam \top/processor/sha_core/hash_out_88_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_87_s0  (
	.D(\top/processor/sha_core/h5 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [87])
);
defparam \top/processor/sha_core/hash_out_87_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_86_s0  (
	.D(\top/processor/sha_core/h5 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [86])
);
defparam \top/processor/sha_core/hash_out_86_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_85_s0  (
	.D(\top/processor/sha_core/h5 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [85])
);
defparam \top/processor/sha_core/hash_out_85_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_84_s0  (
	.D(\top/processor/sha_core/h5 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [84])
);
defparam \top/processor/sha_core/hash_out_84_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_83_s0  (
	.D(\top/processor/sha_core/h5 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [83])
);
defparam \top/processor/sha_core/hash_out_83_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_82_s0  (
	.D(\top/processor/sha_core/h5 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [82])
);
defparam \top/processor/sha_core/hash_out_82_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_81_s0  (
	.D(\top/processor/sha_core/h5 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [81])
);
defparam \top/processor/sha_core/hash_out_81_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_80_s0  (
	.D(\top/processor/sha_core/h5 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [80])
);
defparam \top/processor/sha_core/hash_out_80_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_79_s0  (
	.D(\top/processor/sha_core/h5 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [79])
);
defparam \top/processor/sha_core/hash_out_79_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_78_s0  (
	.D(\top/processor/sha_core/h5 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [78])
);
defparam \top/processor/sha_core/hash_out_78_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_77_s0  (
	.D(\top/processor/sha_core/h5 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [77])
);
defparam \top/processor/sha_core/hash_out_77_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_76_s0  (
	.D(\top/processor/sha_core/h5 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [76])
);
defparam \top/processor/sha_core/hash_out_76_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_75_s0  (
	.D(\top/processor/sha_core/h5 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [75])
);
defparam \top/processor/sha_core/hash_out_75_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_74_s0  (
	.D(\top/processor/sha_core/h5 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [74])
);
defparam \top/processor/sha_core/hash_out_74_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_73_s0  (
	.D(\top/processor/sha_core/h5 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [73])
);
defparam \top/processor/sha_core/hash_out_73_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_72_s0  (
	.D(\top/processor/sha_core/h5 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [72])
);
defparam \top/processor/sha_core/hash_out_72_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_71_s0  (
	.D(\top/processor/sha_core/h5 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [71])
);
defparam \top/processor/sha_core/hash_out_71_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_70_s0  (
	.D(\top/processor/sha_core/h5 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [70])
);
defparam \top/processor/sha_core/hash_out_70_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_69_s0  (
	.D(\top/processor/sha_core/h5 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [69])
);
defparam \top/processor/sha_core/hash_out_69_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_68_s0  (
	.D(\top/processor/sha_core/h5 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [68])
);
defparam \top/processor/sha_core/hash_out_68_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_67_s0  (
	.D(\top/processor/sha_core/h5 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [67])
);
defparam \top/processor/sha_core/hash_out_67_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_66_s0  (
	.D(\top/processor/sha_core/h5 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [66])
);
defparam \top/processor/sha_core/hash_out_66_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_65_s0  (
	.D(\top/processor/sha_core/h5 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [65])
);
defparam \top/processor/sha_core/hash_out_65_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_64_s0  (
	.D(\top/processor/sha_core/h5 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [64])
);
defparam \top/processor/sha_core/hash_out_64_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_63_s0  (
	.D(\top/processor/sha_core/h6 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [63])
);
defparam \top/processor/sha_core/hash_out_63_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_62_s0  (
	.D(\top/processor/sha_core/h6 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [62])
);
defparam \top/processor/sha_core/hash_out_62_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_61_s0  (
	.D(\top/processor/sha_core/h6 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [61])
);
defparam \top/processor/sha_core/hash_out_61_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_60_s0  (
	.D(\top/processor/sha_core/h6 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [60])
);
defparam \top/processor/sha_core/hash_out_60_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_59_s0  (
	.D(\top/processor/sha_core/h6 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [59])
);
defparam \top/processor/sha_core/hash_out_59_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_58_s0  (
	.D(\top/processor/sha_core/h6 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [58])
);
defparam \top/processor/sha_core/hash_out_58_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_57_s0  (
	.D(\top/processor/sha_core/h6 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [57])
);
defparam \top/processor/sha_core/hash_out_57_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_56_s0  (
	.D(\top/processor/sha_core/h6 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [56])
);
defparam \top/processor/sha_core/hash_out_56_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_55_s0  (
	.D(\top/processor/sha_core/h6 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [55])
);
defparam \top/processor/sha_core/hash_out_55_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_54_s0  (
	.D(\top/processor/sha_core/h6 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [54])
);
defparam \top/processor/sha_core/hash_out_54_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_53_s0  (
	.D(\top/processor/sha_core/h6 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [53])
);
defparam \top/processor/sha_core/hash_out_53_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_52_s0  (
	.D(\top/processor/sha_core/h6 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [52])
);
defparam \top/processor/sha_core/hash_out_52_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_51_s0  (
	.D(\top/processor/sha_core/h6 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [51])
);
defparam \top/processor/sha_core/hash_out_51_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_50_s0  (
	.D(\top/processor/sha_core/h6 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [50])
);
defparam \top/processor/sha_core/hash_out_50_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_49_s0  (
	.D(\top/processor/sha_core/h6 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [49])
);
defparam \top/processor/sha_core/hash_out_49_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_48_s0  (
	.D(\top/processor/sha_core/h6 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [48])
);
defparam \top/processor/sha_core/hash_out_48_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_47_s0  (
	.D(\top/processor/sha_core/h6 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [47])
);
defparam \top/processor/sha_core/hash_out_47_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_46_s0  (
	.D(\top/processor/sha_core/h6 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [46])
);
defparam \top/processor/sha_core/hash_out_46_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_45_s0  (
	.D(\top/processor/sha_core/h6 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [45])
);
defparam \top/processor/sha_core/hash_out_45_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_44_s0  (
	.D(\top/processor/sha_core/h6 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [44])
);
defparam \top/processor/sha_core/hash_out_44_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_43_s0  (
	.D(\top/processor/sha_core/h6 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [43])
);
defparam \top/processor/sha_core/hash_out_43_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_42_s0  (
	.D(\top/processor/sha_core/h6 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [42])
);
defparam \top/processor/sha_core/hash_out_42_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_41_s0  (
	.D(\top/processor/sha_core/h6 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [41])
);
defparam \top/processor/sha_core/hash_out_41_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_40_s0  (
	.D(\top/processor/sha_core/h6 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [40])
);
defparam \top/processor/sha_core/hash_out_40_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_39_s0  (
	.D(\top/processor/sha_core/h6 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [39])
);
defparam \top/processor/sha_core/hash_out_39_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_38_s0  (
	.D(\top/processor/sha_core/h6 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [38])
);
defparam \top/processor/sha_core/hash_out_38_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_37_s0  (
	.D(\top/processor/sha_core/h6 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [37])
);
defparam \top/processor/sha_core/hash_out_37_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_36_s0  (
	.D(\top/processor/sha_core/h6 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [36])
);
defparam \top/processor/sha_core/hash_out_36_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_35_s0  (
	.D(\top/processor/sha_core/h6 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [35])
);
defparam \top/processor/sha_core/hash_out_35_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_34_s0  (
	.D(\top/processor/sha_core/h6 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [34])
);
defparam \top/processor/sha_core/hash_out_34_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_33_s0  (
	.D(\top/processor/sha_core/h6 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [33])
);
defparam \top/processor/sha_core/hash_out_33_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_32_s0  (
	.D(\top/processor/sha_core/h6 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [32])
);
defparam \top/processor/sha_core/hash_out_32_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_31_s0  (
	.D(\top/processor/sha_core/h7 [31]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [31])
);
defparam \top/processor/sha_core/hash_out_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_30_s0  (
	.D(\top/processor/sha_core/h7 [30]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [30])
);
defparam \top/processor/sha_core/hash_out_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_29_s0  (
	.D(\top/processor/sha_core/h7 [29]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [29])
);
defparam \top/processor/sha_core/hash_out_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_28_s0  (
	.D(\top/processor/sha_core/h7 [28]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [28])
);
defparam \top/processor/sha_core/hash_out_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_27_s0  (
	.D(\top/processor/sha_core/h7 [27]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [27])
);
defparam \top/processor/sha_core/hash_out_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_26_s0  (
	.D(\top/processor/sha_core/h7 [26]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [26])
);
defparam \top/processor/sha_core/hash_out_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_25_s0  (
	.D(\top/processor/sha_core/h7 [25]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [25])
);
defparam \top/processor/sha_core/hash_out_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_24_s0  (
	.D(\top/processor/sha_core/h7 [24]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [24])
);
defparam \top/processor/sha_core/hash_out_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_23_s0  (
	.D(\top/processor/sha_core/h7 [23]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [23])
);
defparam \top/processor/sha_core/hash_out_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_22_s0  (
	.D(\top/processor/sha_core/h7 [22]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [22])
);
defparam \top/processor/sha_core/hash_out_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_21_s0  (
	.D(\top/processor/sha_core/h7 [21]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [21])
);
defparam \top/processor/sha_core/hash_out_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_20_s0  (
	.D(\top/processor/sha_core/h7 [20]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [20])
);
defparam \top/processor/sha_core/hash_out_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_19_s0  (
	.D(\top/processor/sha_core/h7 [19]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [19])
);
defparam \top/processor/sha_core/hash_out_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_18_s0  (
	.D(\top/processor/sha_core/h7 [18]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [18])
);
defparam \top/processor/sha_core/hash_out_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_17_s0  (
	.D(\top/processor/sha_core/h7 [17]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [17])
);
defparam \top/processor/sha_core/hash_out_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_16_s0  (
	.D(\top/processor/sha_core/h7 [16]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [16])
);
defparam \top/processor/sha_core/hash_out_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_15_s0  (
	.D(\top/processor/sha_core/h7 [15]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [15])
);
defparam \top/processor/sha_core/hash_out_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_14_s0  (
	.D(\top/processor/sha_core/h7 [14]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [14])
);
defparam \top/processor/sha_core/hash_out_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_13_s0  (
	.D(\top/processor/sha_core/h7 [13]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [13])
);
defparam \top/processor/sha_core/hash_out_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_12_s0  (
	.D(\top/processor/sha_core/h7 [12]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [12])
);
defparam \top/processor/sha_core/hash_out_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_11_s0  (
	.D(\top/processor/sha_core/h7 [11]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [11])
);
defparam \top/processor/sha_core/hash_out_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_10_s0  (
	.D(\top/processor/sha_core/h7 [10]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [10])
);
defparam \top/processor/sha_core/hash_out_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_9_s0  (
	.D(\top/processor/sha_core/h7 [9]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [9])
);
defparam \top/processor/sha_core/hash_out_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_8_s0  (
	.D(\top/processor/sha_core/h7 [8]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [8])
);
defparam \top/processor/sha_core/hash_out_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_7_s0  (
	.D(\top/processor/sha_core/h7 [7]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [7])
);
defparam \top/processor/sha_core/hash_out_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_6_s0  (
	.D(\top/processor/sha_core/h7 [6]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [6])
);
defparam \top/processor/sha_core/hash_out_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_5_s0  (
	.D(\top/processor/sha_core/h7 [5]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [5])
);
defparam \top/processor/sha_core/hash_out_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_4_s0  (
	.D(\top/processor/sha_core/h7 [4]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [4])
);
defparam \top/processor/sha_core/hash_out_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_3_s0  (
	.D(\top/processor/sha_core/h7 [3]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [3])
);
defparam \top/processor/sha_core/hash_out_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_2_s0  (
	.D(\top/processor/sha_core/h7 [2]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [2])
);
defparam \top/processor/sha_core/hash_out_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_1_s0  (
	.D(\top/processor/sha_core/h7 [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [1])
);
defparam \top/processor/sha_core/hash_out_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/hash_out_0_s0  (
	.D(\top/processor/sha_core/h7 [0]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11613_8 ),
	.CLEAR(rst),
	.Q(\top/processor/core_hash_out [0])
);
defparam \top/processor/sha_core/hash_out_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_6_s0  (
	.D(\top/processor/sha_core/n14439_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [6])
);
defparam \top/processor/sha_core/msg_idx_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_5_s0  (
	.D(\top/processor/sha_core/n14440_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [5])
);
defparam \top/processor/sha_core/msg_idx_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_4_s0  (
	.D(\top/processor/sha_core/n14441_12 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [4])
);
defparam \top/processor/sha_core/msg_idx_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_3_s0  (
	.D(\top/processor/sha_core/n14442_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [3])
);
defparam \top/processor/sha_core/msg_idx_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_2_s0  (
	.D(\top/processor/sha_core/n14443_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [2])
);
defparam \top/processor/sha_core/msg_idx_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_1_s0  (
	.D(\top/processor/sha_core/n14444_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [1])
);
defparam \top/processor/sha_core/msg_idx_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/msg_idx_0_s0  (
	.D(\top/processor/sha_core/n14445_10 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/msg_idx_6_7 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/msg_idx [0])
);
defparam \top/processor/sha_core/msg_idx_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [31])
);
defparam \top/processor/sha_core/w[0]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [30])
);
defparam \top/processor/sha_core/w[0]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [29])
);
defparam \top/processor/sha_core/w[0]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [28])
);
defparam \top/processor/sha_core/w[0]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [27])
);
defparam \top/processor/sha_core/w[0]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [26])
);
defparam \top/processor/sha_core/w[0]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [25])
);
defparam \top/processor/sha_core/w[0]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [24])
);
defparam \top/processor/sha_core/w[0]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [23])
);
defparam \top/processor/sha_core/w[0]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [22])
);
defparam \top/processor/sha_core/w[0]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [21])
);
defparam \top/processor/sha_core/w[0]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [20])
);
defparam \top/processor/sha_core/w[0]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [19])
);
defparam \top/processor/sha_core/w[0]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [18])
);
defparam \top/processor/sha_core/w[0]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [17])
);
defparam \top/processor/sha_core/w[0]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [16])
);
defparam \top/processor/sha_core/w[0]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [15])
);
defparam \top/processor/sha_core/w[0]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [14])
);
defparam \top/processor/sha_core/w[0]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [13])
);
defparam \top/processor/sha_core/w[0]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [12])
);
defparam \top/processor/sha_core/w[0]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [11])
);
defparam \top/processor/sha_core/w[0]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [10])
);
defparam \top/processor/sha_core/w[0]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [9])
);
defparam \top/processor/sha_core/w[0]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [8])
);
defparam \top/processor/sha_core/w[0]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [7])
);
defparam \top/processor/sha_core/w[0]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [6])
);
defparam \top/processor/sha_core/w[0]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [5])
);
defparam \top/processor/sha_core/w[0]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [4])
);
defparam \top/processor/sha_core/w[0]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [3])
);
defparam \top/processor/sha_core/w[0]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [2])
);
defparam \top/processor/sha_core/w[0]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [1])
);
defparam \top/processor/sha_core/w[0]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[0]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[0]_31_12 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[0] [0])
);
defparam \top/processor/sha_core/w[0]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [31])
);
defparam \top/processor/sha_core/w[1]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [30])
);
defparam \top/processor/sha_core/w[1]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [29])
);
defparam \top/processor/sha_core/w[1]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [28])
);
defparam \top/processor/sha_core/w[1]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [27])
);
defparam \top/processor/sha_core/w[1]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [26])
);
defparam \top/processor/sha_core/w[1]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [25])
);
defparam \top/processor/sha_core/w[1]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [24])
);
defparam \top/processor/sha_core/w[1]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [23])
);
defparam \top/processor/sha_core/w[1]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [22])
);
defparam \top/processor/sha_core/w[1]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [21])
);
defparam \top/processor/sha_core/w[1]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [20])
);
defparam \top/processor/sha_core/w[1]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [19])
);
defparam \top/processor/sha_core/w[1]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [18])
);
defparam \top/processor/sha_core/w[1]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [17])
);
defparam \top/processor/sha_core/w[1]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [16])
);
defparam \top/processor/sha_core/w[1]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [15])
);
defparam \top/processor/sha_core/w[1]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [14])
);
defparam \top/processor/sha_core/w[1]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [13])
);
defparam \top/processor/sha_core/w[1]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [12])
);
defparam \top/processor/sha_core/w[1]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [11])
);
defparam \top/processor/sha_core/w[1]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [10])
);
defparam \top/processor/sha_core/w[1]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [9])
);
defparam \top/processor/sha_core/w[1]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [8])
);
defparam \top/processor/sha_core/w[1]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [7])
);
defparam \top/processor/sha_core/w[1]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [6])
);
defparam \top/processor/sha_core/w[1]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [5])
);
defparam \top/processor/sha_core/w[1]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [4])
);
defparam \top/processor/sha_core/w[1]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [3])
);
defparam \top/processor/sha_core/w[1]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [2])
);
defparam \top/processor/sha_core/w[1]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [1])
);
defparam \top/processor/sha_core/w[1]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[1]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[1]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[1] [0])
);
defparam \top/processor/sha_core/w[1]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [31])
);
defparam \top/processor/sha_core/w[2]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [30])
);
defparam \top/processor/sha_core/w[2]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [29])
);
defparam \top/processor/sha_core/w[2]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [28])
);
defparam \top/processor/sha_core/w[2]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [27])
);
defparam \top/processor/sha_core/w[2]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [26])
);
defparam \top/processor/sha_core/w[2]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [25])
);
defparam \top/processor/sha_core/w[2]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [24])
);
defparam \top/processor/sha_core/w[2]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [23])
);
defparam \top/processor/sha_core/w[2]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [22])
);
defparam \top/processor/sha_core/w[2]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [21])
);
defparam \top/processor/sha_core/w[2]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [20])
);
defparam \top/processor/sha_core/w[2]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [19])
);
defparam \top/processor/sha_core/w[2]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [18])
);
defparam \top/processor/sha_core/w[2]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [17])
);
defparam \top/processor/sha_core/w[2]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [16])
);
defparam \top/processor/sha_core/w[2]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [15])
);
defparam \top/processor/sha_core/w[2]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [14])
);
defparam \top/processor/sha_core/w[2]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [13])
);
defparam \top/processor/sha_core/w[2]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [12])
);
defparam \top/processor/sha_core/w[2]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [11])
);
defparam \top/processor/sha_core/w[2]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [10])
);
defparam \top/processor/sha_core/w[2]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [9])
);
defparam \top/processor/sha_core/w[2]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [8])
);
defparam \top/processor/sha_core/w[2]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [7])
);
defparam \top/processor/sha_core/w[2]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [6])
);
defparam \top/processor/sha_core/w[2]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [5])
);
defparam \top/processor/sha_core/w[2]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [4])
);
defparam \top/processor/sha_core/w[2]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [3])
);
defparam \top/processor/sha_core/w[2]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [2])
);
defparam \top/processor/sha_core/w[2]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [1])
);
defparam \top/processor/sha_core/w[2]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[2]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[2]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[2] [0])
);
defparam \top/processor/sha_core/w[2]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [31])
);
defparam \top/processor/sha_core/w[3]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [30])
);
defparam \top/processor/sha_core/w[3]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [29])
);
defparam \top/processor/sha_core/w[3]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [28])
);
defparam \top/processor/sha_core/w[3]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [27])
);
defparam \top/processor/sha_core/w[3]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [26])
);
defparam \top/processor/sha_core/w[3]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [25])
);
defparam \top/processor/sha_core/w[3]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [24])
);
defparam \top/processor/sha_core/w[3]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [23])
);
defparam \top/processor/sha_core/w[3]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [22])
);
defparam \top/processor/sha_core/w[3]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [21])
);
defparam \top/processor/sha_core/w[3]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [20])
);
defparam \top/processor/sha_core/w[3]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [19])
);
defparam \top/processor/sha_core/w[3]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [18])
);
defparam \top/processor/sha_core/w[3]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [17])
);
defparam \top/processor/sha_core/w[3]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [16])
);
defparam \top/processor/sha_core/w[3]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [15])
);
defparam \top/processor/sha_core/w[3]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [14])
);
defparam \top/processor/sha_core/w[3]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [13])
);
defparam \top/processor/sha_core/w[3]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [12])
);
defparam \top/processor/sha_core/w[3]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [11])
);
defparam \top/processor/sha_core/w[3]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [10])
);
defparam \top/processor/sha_core/w[3]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [9])
);
defparam \top/processor/sha_core/w[3]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [8])
);
defparam \top/processor/sha_core/w[3]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [7])
);
defparam \top/processor/sha_core/w[3]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [6])
);
defparam \top/processor/sha_core/w[3]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [5])
);
defparam \top/processor/sha_core/w[3]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [4])
);
defparam \top/processor/sha_core/w[3]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [3])
);
defparam \top/processor/sha_core/w[3]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [2])
);
defparam \top/processor/sha_core/w[3]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [1])
);
defparam \top/processor/sha_core/w[3]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[3]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[3]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[3] [0])
);
defparam \top/processor/sha_core/w[3]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [31])
);
defparam \top/processor/sha_core/w[4]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [30])
);
defparam \top/processor/sha_core/w[4]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [29])
);
defparam \top/processor/sha_core/w[4]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [28])
);
defparam \top/processor/sha_core/w[4]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [27])
);
defparam \top/processor/sha_core/w[4]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [26])
);
defparam \top/processor/sha_core/w[4]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [25])
);
defparam \top/processor/sha_core/w[4]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [24])
);
defparam \top/processor/sha_core/w[4]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [23])
);
defparam \top/processor/sha_core/w[4]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [22])
);
defparam \top/processor/sha_core/w[4]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [21])
);
defparam \top/processor/sha_core/w[4]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [20])
);
defparam \top/processor/sha_core/w[4]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [19])
);
defparam \top/processor/sha_core/w[4]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [18])
);
defparam \top/processor/sha_core/w[4]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [17])
);
defparam \top/processor/sha_core/w[4]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [16])
);
defparam \top/processor/sha_core/w[4]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [15])
);
defparam \top/processor/sha_core/w[4]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [14])
);
defparam \top/processor/sha_core/w[4]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [13])
);
defparam \top/processor/sha_core/w[4]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [12])
);
defparam \top/processor/sha_core/w[4]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [11])
);
defparam \top/processor/sha_core/w[4]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [10])
);
defparam \top/processor/sha_core/w[4]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [9])
);
defparam \top/processor/sha_core/w[4]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [8])
);
defparam \top/processor/sha_core/w[4]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [7])
);
defparam \top/processor/sha_core/w[4]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [6])
);
defparam \top/processor/sha_core/w[4]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [5])
);
defparam \top/processor/sha_core/w[4]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [4])
);
defparam \top/processor/sha_core/w[4]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [3])
);
defparam \top/processor/sha_core/w[4]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [2])
);
defparam \top/processor/sha_core/w[4]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [1])
);
defparam \top/processor/sha_core/w[4]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[4]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[4]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[4] [0])
);
defparam \top/processor/sha_core/w[4]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [31])
);
defparam \top/processor/sha_core/w[5]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [30])
);
defparam \top/processor/sha_core/w[5]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [29])
);
defparam \top/processor/sha_core/w[5]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [28])
);
defparam \top/processor/sha_core/w[5]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [27])
);
defparam \top/processor/sha_core/w[5]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [26])
);
defparam \top/processor/sha_core/w[5]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [25])
);
defparam \top/processor/sha_core/w[5]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [24])
);
defparam \top/processor/sha_core/w[5]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [23])
);
defparam \top/processor/sha_core/w[5]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [22])
);
defparam \top/processor/sha_core/w[5]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [21])
);
defparam \top/processor/sha_core/w[5]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [20])
);
defparam \top/processor/sha_core/w[5]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [19])
);
defparam \top/processor/sha_core/w[5]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [18])
);
defparam \top/processor/sha_core/w[5]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [17])
);
defparam \top/processor/sha_core/w[5]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [16])
);
defparam \top/processor/sha_core/w[5]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [15])
);
defparam \top/processor/sha_core/w[5]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [14])
);
defparam \top/processor/sha_core/w[5]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [13])
);
defparam \top/processor/sha_core/w[5]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [12])
);
defparam \top/processor/sha_core/w[5]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [11])
);
defparam \top/processor/sha_core/w[5]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [10])
);
defparam \top/processor/sha_core/w[5]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [9])
);
defparam \top/processor/sha_core/w[5]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [8])
);
defparam \top/processor/sha_core/w[5]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [7])
);
defparam \top/processor/sha_core/w[5]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [6])
);
defparam \top/processor/sha_core/w[5]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [5])
);
defparam \top/processor/sha_core/w[5]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [4])
);
defparam \top/processor/sha_core/w[5]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [3])
);
defparam \top/processor/sha_core/w[5]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [2])
);
defparam \top/processor/sha_core/w[5]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [1])
);
defparam \top/processor/sha_core/w[5]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[5]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[5]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[5] [0])
);
defparam \top/processor/sha_core/w[5]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [31])
);
defparam \top/processor/sha_core/w[6]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [30])
);
defparam \top/processor/sha_core/w[6]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [29])
);
defparam \top/processor/sha_core/w[6]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [28])
);
defparam \top/processor/sha_core/w[6]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [27])
);
defparam \top/processor/sha_core/w[6]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [26])
);
defparam \top/processor/sha_core/w[6]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [25])
);
defparam \top/processor/sha_core/w[6]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [24])
);
defparam \top/processor/sha_core/w[6]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [23])
);
defparam \top/processor/sha_core/w[6]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [22])
);
defparam \top/processor/sha_core/w[6]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [21])
);
defparam \top/processor/sha_core/w[6]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [20])
);
defparam \top/processor/sha_core/w[6]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [19])
);
defparam \top/processor/sha_core/w[6]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [18])
);
defparam \top/processor/sha_core/w[6]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [17])
);
defparam \top/processor/sha_core/w[6]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [16])
);
defparam \top/processor/sha_core/w[6]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [15])
);
defparam \top/processor/sha_core/w[6]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [14])
);
defparam \top/processor/sha_core/w[6]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [13])
);
defparam \top/processor/sha_core/w[6]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [12])
);
defparam \top/processor/sha_core/w[6]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [11])
);
defparam \top/processor/sha_core/w[6]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [10])
);
defparam \top/processor/sha_core/w[6]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [9])
);
defparam \top/processor/sha_core/w[6]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [8])
);
defparam \top/processor/sha_core/w[6]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [7])
);
defparam \top/processor/sha_core/w[6]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [6])
);
defparam \top/processor/sha_core/w[6]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [5])
);
defparam \top/processor/sha_core/w[6]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [4])
);
defparam \top/processor/sha_core/w[6]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [3])
);
defparam \top/processor/sha_core/w[6]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [2])
);
defparam \top/processor/sha_core/w[6]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [1])
);
defparam \top/processor/sha_core/w[6]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[6]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[6]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[6] [0])
);
defparam \top/processor/sha_core/w[6]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [31])
);
defparam \top/processor/sha_core/w[7]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [30])
);
defparam \top/processor/sha_core/w[7]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [29])
);
defparam \top/processor/sha_core/w[7]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [28])
);
defparam \top/processor/sha_core/w[7]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [27])
);
defparam \top/processor/sha_core/w[7]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [26])
);
defparam \top/processor/sha_core/w[7]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [25])
);
defparam \top/processor/sha_core/w[7]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [24])
);
defparam \top/processor/sha_core/w[7]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [23])
);
defparam \top/processor/sha_core/w[7]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [22])
);
defparam \top/processor/sha_core/w[7]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [21])
);
defparam \top/processor/sha_core/w[7]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [20])
);
defparam \top/processor/sha_core/w[7]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [19])
);
defparam \top/processor/sha_core/w[7]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [18])
);
defparam \top/processor/sha_core/w[7]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [17])
);
defparam \top/processor/sha_core/w[7]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [16])
);
defparam \top/processor/sha_core/w[7]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [15])
);
defparam \top/processor/sha_core/w[7]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [14])
);
defparam \top/processor/sha_core/w[7]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [13])
);
defparam \top/processor/sha_core/w[7]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [12])
);
defparam \top/processor/sha_core/w[7]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [11])
);
defparam \top/processor/sha_core/w[7]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [10])
);
defparam \top/processor/sha_core/w[7]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [9])
);
defparam \top/processor/sha_core/w[7]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [8])
);
defparam \top/processor/sha_core/w[7]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [7])
);
defparam \top/processor/sha_core/w[7]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [6])
);
defparam \top/processor/sha_core/w[7]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [5])
);
defparam \top/processor/sha_core/w[7]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [4])
);
defparam \top/processor/sha_core/w[7]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [3])
);
defparam \top/processor/sha_core/w[7]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [2])
);
defparam \top/processor/sha_core/w[7]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [1])
);
defparam \top/processor/sha_core/w[7]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[7]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[7]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[7] [0])
);
defparam \top/processor/sha_core/w[7]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [31])
);
defparam \top/processor/sha_core/w[8]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [30])
);
defparam \top/processor/sha_core/w[8]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [29])
);
defparam \top/processor/sha_core/w[8]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [28])
);
defparam \top/processor/sha_core/w[8]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [27])
);
defparam \top/processor/sha_core/w[8]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [26])
);
defparam \top/processor/sha_core/w[8]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [25])
);
defparam \top/processor/sha_core/w[8]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [24])
);
defparam \top/processor/sha_core/w[8]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [23])
);
defparam \top/processor/sha_core/w[8]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [22])
);
defparam \top/processor/sha_core/w[8]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [21])
);
defparam \top/processor/sha_core/w[8]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [20])
);
defparam \top/processor/sha_core/w[8]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [19])
);
defparam \top/processor/sha_core/w[8]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [18])
);
defparam \top/processor/sha_core/w[8]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [17])
);
defparam \top/processor/sha_core/w[8]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [16])
);
defparam \top/processor/sha_core/w[8]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [15])
);
defparam \top/processor/sha_core/w[8]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [14])
);
defparam \top/processor/sha_core/w[8]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [13])
);
defparam \top/processor/sha_core/w[8]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [12])
);
defparam \top/processor/sha_core/w[8]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [11])
);
defparam \top/processor/sha_core/w[8]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [10])
);
defparam \top/processor/sha_core/w[8]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [9])
);
defparam \top/processor/sha_core/w[8]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [8])
);
defparam \top/processor/sha_core/w[8]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [7])
);
defparam \top/processor/sha_core/w[8]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [6])
);
defparam \top/processor/sha_core/w[8]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [5])
);
defparam \top/processor/sha_core/w[8]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [4])
);
defparam \top/processor/sha_core/w[8]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [3])
);
defparam \top/processor/sha_core/w[8]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [2])
);
defparam \top/processor/sha_core/w[8]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [1])
);
defparam \top/processor/sha_core/w[8]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[8]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[8]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[8] [0])
);
defparam \top/processor/sha_core/w[8]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [31])
);
defparam \top/processor/sha_core/w[9]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [30])
);
defparam \top/processor/sha_core/w[9]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [29])
);
defparam \top/processor/sha_core/w[9]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [28])
);
defparam \top/processor/sha_core/w[9]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [27])
);
defparam \top/processor/sha_core/w[9]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [26])
);
defparam \top/processor/sha_core/w[9]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [25])
);
defparam \top/processor/sha_core/w[9]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [24])
);
defparam \top/processor/sha_core/w[9]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [23])
);
defparam \top/processor/sha_core/w[9]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [22])
);
defparam \top/processor/sha_core/w[9]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [21])
);
defparam \top/processor/sha_core/w[9]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [20])
);
defparam \top/processor/sha_core/w[9]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [19])
);
defparam \top/processor/sha_core/w[9]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [18])
);
defparam \top/processor/sha_core/w[9]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [17])
);
defparam \top/processor/sha_core/w[9]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [16])
);
defparam \top/processor/sha_core/w[9]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [15])
);
defparam \top/processor/sha_core/w[9]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [14])
);
defparam \top/processor/sha_core/w[9]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [13])
);
defparam \top/processor/sha_core/w[9]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [12])
);
defparam \top/processor/sha_core/w[9]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [11])
);
defparam \top/processor/sha_core/w[9]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [10])
);
defparam \top/processor/sha_core/w[9]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [9])
);
defparam \top/processor/sha_core/w[9]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [8])
);
defparam \top/processor/sha_core/w[9]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [7])
);
defparam \top/processor/sha_core/w[9]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [6])
);
defparam \top/processor/sha_core/w[9]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [5])
);
defparam \top/processor/sha_core/w[9]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [4])
);
defparam \top/processor/sha_core/w[9]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [3])
);
defparam \top/processor/sha_core/w[9]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [2])
);
defparam \top/processor/sha_core/w[9]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [1])
);
defparam \top/processor/sha_core/w[9]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[9]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[9]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[9] [0])
);
defparam \top/processor/sha_core/w[9]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [31])
);
defparam \top/processor/sha_core/w[10]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [30])
);
defparam \top/processor/sha_core/w[10]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [29])
);
defparam \top/processor/sha_core/w[10]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [28])
);
defparam \top/processor/sha_core/w[10]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [27])
);
defparam \top/processor/sha_core/w[10]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [26])
);
defparam \top/processor/sha_core/w[10]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [25])
);
defparam \top/processor/sha_core/w[10]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [24])
);
defparam \top/processor/sha_core/w[10]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [23])
);
defparam \top/processor/sha_core/w[10]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [22])
);
defparam \top/processor/sha_core/w[10]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [21])
);
defparam \top/processor/sha_core/w[10]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [20])
);
defparam \top/processor/sha_core/w[10]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [19])
);
defparam \top/processor/sha_core/w[10]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [18])
);
defparam \top/processor/sha_core/w[10]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [17])
);
defparam \top/processor/sha_core/w[10]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [16])
);
defparam \top/processor/sha_core/w[10]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [15])
);
defparam \top/processor/sha_core/w[10]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [14])
);
defparam \top/processor/sha_core/w[10]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [13])
);
defparam \top/processor/sha_core/w[10]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [12])
);
defparam \top/processor/sha_core/w[10]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [11])
);
defparam \top/processor/sha_core/w[10]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [10])
);
defparam \top/processor/sha_core/w[10]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [9])
);
defparam \top/processor/sha_core/w[10]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [8])
);
defparam \top/processor/sha_core/w[10]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [7])
);
defparam \top/processor/sha_core/w[10]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [6])
);
defparam \top/processor/sha_core/w[10]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [5])
);
defparam \top/processor/sha_core/w[10]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [4])
);
defparam \top/processor/sha_core/w[10]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [3])
);
defparam \top/processor/sha_core/w[10]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [2])
);
defparam \top/processor/sha_core/w[10]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [1])
);
defparam \top/processor/sha_core/w[10]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[10]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[10]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[10] [0])
);
defparam \top/processor/sha_core/w[10]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [31])
);
defparam \top/processor/sha_core/w[11]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [30])
);
defparam \top/processor/sha_core/w[11]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [29])
);
defparam \top/processor/sha_core/w[11]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [28])
);
defparam \top/processor/sha_core/w[11]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [27])
);
defparam \top/processor/sha_core/w[11]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [26])
);
defparam \top/processor/sha_core/w[11]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [25])
);
defparam \top/processor/sha_core/w[11]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [24])
);
defparam \top/processor/sha_core/w[11]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [23])
);
defparam \top/processor/sha_core/w[11]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [22])
);
defparam \top/processor/sha_core/w[11]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [21])
);
defparam \top/processor/sha_core/w[11]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [20])
);
defparam \top/processor/sha_core/w[11]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [19])
);
defparam \top/processor/sha_core/w[11]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [18])
);
defparam \top/processor/sha_core/w[11]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [17])
);
defparam \top/processor/sha_core/w[11]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [16])
);
defparam \top/processor/sha_core/w[11]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [15])
);
defparam \top/processor/sha_core/w[11]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [14])
);
defparam \top/processor/sha_core/w[11]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [13])
);
defparam \top/processor/sha_core/w[11]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [12])
);
defparam \top/processor/sha_core/w[11]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [11])
);
defparam \top/processor/sha_core/w[11]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [10])
);
defparam \top/processor/sha_core/w[11]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [9])
);
defparam \top/processor/sha_core/w[11]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [8])
);
defparam \top/processor/sha_core/w[11]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [7])
);
defparam \top/processor/sha_core/w[11]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [6])
);
defparam \top/processor/sha_core/w[11]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [5])
);
defparam \top/processor/sha_core/w[11]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [4])
);
defparam \top/processor/sha_core/w[11]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [3])
);
defparam \top/processor/sha_core/w[11]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [2])
);
defparam \top/processor/sha_core/w[11]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [1])
);
defparam \top/processor/sha_core/w[11]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[11]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[11]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[11] [0])
);
defparam \top/processor/sha_core/w[11]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [31])
);
defparam \top/processor/sha_core/w[12]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [30])
);
defparam \top/processor/sha_core/w[12]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [29])
);
defparam \top/processor/sha_core/w[12]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [28])
);
defparam \top/processor/sha_core/w[12]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [27])
);
defparam \top/processor/sha_core/w[12]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [26])
);
defparam \top/processor/sha_core/w[12]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [25])
);
defparam \top/processor/sha_core/w[12]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [24])
);
defparam \top/processor/sha_core/w[12]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [23])
);
defparam \top/processor/sha_core/w[12]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [22])
);
defparam \top/processor/sha_core/w[12]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [21])
);
defparam \top/processor/sha_core/w[12]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [20])
);
defparam \top/processor/sha_core/w[12]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [19])
);
defparam \top/processor/sha_core/w[12]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [18])
);
defparam \top/processor/sha_core/w[12]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [17])
);
defparam \top/processor/sha_core/w[12]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [16])
);
defparam \top/processor/sha_core/w[12]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [15])
);
defparam \top/processor/sha_core/w[12]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [14])
);
defparam \top/processor/sha_core/w[12]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [13])
);
defparam \top/processor/sha_core/w[12]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [12])
);
defparam \top/processor/sha_core/w[12]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [11])
);
defparam \top/processor/sha_core/w[12]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [10])
);
defparam \top/processor/sha_core/w[12]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [9])
);
defparam \top/processor/sha_core/w[12]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [8])
);
defparam \top/processor/sha_core/w[12]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [7])
);
defparam \top/processor/sha_core/w[12]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [6])
);
defparam \top/processor/sha_core/w[12]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [5])
);
defparam \top/processor/sha_core/w[12]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [4])
);
defparam \top/processor/sha_core/w[12]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [3])
);
defparam \top/processor/sha_core/w[12]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [2])
);
defparam \top/processor/sha_core/w[12]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [1])
);
defparam \top/processor/sha_core/w[12]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[12]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[12]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[12] [0])
);
defparam \top/processor/sha_core/w[12]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [31])
);
defparam \top/processor/sha_core/w[13]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [30])
);
defparam \top/processor/sha_core/w[13]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [29])
);
defparam \top/processor/sha_core/w[13]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [28])
);
defparam \top/processor/sha_core/w[13]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [27])
);
defparam \top/processor/sha_core/w[13]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [26])
);
defparam \top/processor/sha_core/w[13]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [25])
);
defparam \top/processor/sha_core/w[13]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [24])
);
defparam \top/processor/sha_core/w[13]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [23])
);
defparam \top/processor/sha_core/w[13]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [22])
);
defparam \top/processor/sha_core/w[13]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [21])
);
defparam \top/processor/sha_core/w[13]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [20])
);
defparam \top/processor/sha_core/w[13]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [19])
);
defparam \top/processor/sha_core/w[13]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [18])
);
defparam \top/processor/sha_core/w[13]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [17])
);
defparam \top/processor/sha_core/w[13]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [16])
);
defparam \top/processor/sha_core/w[13]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [15])
);
defparam \top/processor/sha_core/w[13]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [14])
);
defparam \top/processor/sha_core/w[13]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [13])
);
defparam \top/processor/sha_core/w[13]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [12])
);
defparam \top/processor/sha_core/w[13]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [11])
);
defparam \top/processor/sha_core/w[13]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [10])
);
defparam \top/processor/sha_core/w[13]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [9])
);
defparam \top/processor/sha_core/w[13]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [8])
);
defparam \top/processor/sha_core/w[13]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [7])
);
defparam \top/processor/sha_core/w[13]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [6])
);
defparam \top/processor/sha_core/w[13]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [5])
);
defparam \top/processor/sha_core/w[13]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [4])
);
defparam \top/processor/sha_core/w[13]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [3])
);
defparam \top/processor/sha_core/w[13]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [2])
);
defparam \top/processor/sha_core/w[13]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [1])
);
defparam \top/processor/sha_core/w[13]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[13]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[13]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[13] [0])
);
defparam \top/processor/sha_core/w[13]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [31])
);
defparam \top/processor/sha_core/w[14]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [30])
);
defparam \top/processor/sha_core/w[14]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [29])
);
defparam \top/processor/sha_core/w[14]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [28])
);
defparam \top/processor/sha_core/w[14]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [27])
);
defparam \top/processor/sha_core/w[14]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [26])
);
defparam \top/processor/sha_core/w[14]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [25])
);
defparam \top/processor/sha_core/w[14]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [24])
);
defparam \top/processor/sha_core/w[14]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [23])
);
defparam \top/processor/sha_core/w[14]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [22])
);
defparam \top/processor/sha_core/w[14]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [21])
);
defparam \top/processor/sha_core/w[14]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [20])
);
defparam \top/processor/sha_core/w[14]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [19])
);
defparam \top/processor/sha_core/w[14]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [18])
);
defparam \top/processor/sha_core/w[14]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [17])
);
defparam \top/processor/sha_core/w[14]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [16])
);
defparam \top/processor/sha_core/w[14]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [15])
);
defparam \top/processor/sha_core/w[14]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [14])
);
defparam \top/processor/sha_core/w[14]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [13])
);
defparam \top/processor/sha_core/w[14]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [12])
);
defparam \top/processor/sha_core/w[14]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [11])
);
defparam \top/processor/sha_core/w[14]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [10])
);
defparam \top/processor/sha_core/w[14]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [9])
);
defparam \top/processor/sha_core/w[14]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [8])
);
defparam \top/processor/sha_core/w[14]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [7])
);
defparam \top/processor/sha_core/w[14]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [6])
);
defparam \top/processor/sha_core/w[14]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [5])
);
defparam \top/processor/sha_core/w[14]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [4])
);
defparam \top/processor/sha_core/w[14]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [3])
);
defparam \top/processor/sha_core/w[14]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [2])
);
defparam \top/processor/sha_core/w[14]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [1])
);
defparam \top/processor/sha_core/w[14]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[14]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[14]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[14] [0])
);
defparam \top/processor/sha_core/w[14]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [31])
);
defparam \top/processor/sha_core/w[15]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [30])
);
defparam \top/processor/sha_core/w[15]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [29])
);
defparam \top/processor/sha_core/w[15]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [28])
);
defparam \top/processor/sha_core/w[15]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [27])
);
defparam \top/processor/sha_core/w[15]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [26])
);
defparam \top/processor/sha_core/w[15]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [25])
);
defparam \top/processor/sha_core/w[15]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [24])
);
defparam \top/processor/sha_core/w[15]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [23])
);
defparam \top/processor/sha_core/w[15]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [22])
);
defparam \top/processor/sha_core/w[15]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [21])
);
defparam \top/processor/sha_core/w[15]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [20])
);
defparam \top/processor/sha_core/w[15]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [19])
);
defparam \top/processor/sha_core/w[15]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [18])
);
defparam \top/processor/sha_core/w[15]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [17])
);
defparam \top/processor/sha_core/w[15]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [16])
);
defparam \top/processor/sha_core/w[15]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [15])
);
defparam \top/processor/sha_core/w[15]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [14])
);
defparam \top/processor/sha_core/w[15]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [13])
);
defparam \top/processor/sha_core/w[15]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [12])
);
defparam \top/processor/sha_core/w[15]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [11])
);
defparam \top/processor/sha_core/w[15]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [10])
);
defparam \top/processor/sha_core/w[15]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [9])
);
defparam \top/processor/sha_core/w[15]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [8])
);
defparam \top/processor/sha_core/w[15]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [7])
);
defparam \top/processor/sha_core/w[15]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [6])
);
defparam \top/processor/sha_core/w[15]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [5])
);
defparam \top/processor/sha_core/w[15]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [4])
);
defparam \top/processor/sha_core/w[15]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [3])
);
defparam \top/processor/sha_core/w[15]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [2])
);
defparam \top/processor/sha_core/w[15]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [1])
);
defparam \top/processor/sha_core/w[15]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[15]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[15]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[15] [0])
);
defparam \top/processor/sha_core/w[15]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [31])
);
defparam \top/processor/sha_core/w[16]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [30])
);
defparam \top/processor/sha_core/w[16]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [29])
);
defparam \top/processor/sha_core/w[16]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [28])
);
defparam \top/processor/sha_core/w[16]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [27])
);
defparam \top/processor/sha_core/w[16]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [26])
);
defparam \top/processor/sha_core/w[16]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [25])
);
defparam \top/processor/sha_core/w[16]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [24])
);
defparam \top/processor/sha_core/w[16]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [23])
);
defparam \top/processor/sha_core/w[16]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [22])
);
defparam \top/processor/sha_core/w[16]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [21])
);
defparam \top/processor/sha_core/w[16]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [20])
);
defparam \top/processor/sha_core/w[16]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [19])
);
defparam \top/processor/sha_core/w[16]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [18])
);
defparam \top/processor/sha_core/w[16]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [17])
);
defparam \top/processor/sha_core/w[16]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [16])
);
defparam \top/processor/sha_core/w[16]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [15])
);
defparam \top/processor/sha_core/w[16]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [14])
);
defparam \top/processor/sha_core/w[16]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [13])
);
defparam \top/processor/sha_core/w[16]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [12])
);
defparam \top/processor/sha_core/w[16]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [11])
);
defparam \top/processor/sha_core/w[16]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [10])
);
defparam \top/processor/sha_core/w[16]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [9])
);
defparam \top/processor/sha_core/w[16]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [8])
);
defparam \top/processor/sha_core/w[16]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [7])
);
defparam \top/processor/sha_core/w[16]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [6])
);
defparam \top/processor/sha_core/w[16]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [5])
);
defparam \top/processor/sha_core/w[16]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [4])
);
defparam \top/processor/sha_core/w[16]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [3])
);
defparam \top/processor/sha_core/w[16]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [2])
);
defparam \top/processor/sha_core/w[16]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [1])
);
defparam \top/processor/sha_core/w[16]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[16]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[16]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[16] [0])
);
defparam \top/processor/sha_core/w[16]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [31])
);
defparam \top/processor/sha_core/w[17]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [30])
);
defparam \top/processor/sha_core/w[17]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [29])
);
defparam \top/processor/sha_core/w[17]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [28])
);
defparam \top/processor/sha_core/w[17]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [27])
);
defparam \top/processor/sha_core/w[17]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [26])
);
defparam \top/processor/sha_core/w[17]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [25])
);
defparam \top/processor/sha_core/w[17]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [24])
);
defparam \top/processor/sha_core/w[17]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [23])
);
defparam \top/processor/sha_core/w[17]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [22])
);
defparam \top/processor/sha_core/w[17]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [21])
);
defparam \top/processor/sha_core/w[17]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [20])
);
defparam \top/processor/sha_core/w[17]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [19])
);
defparam \top/processor/sha_core/w[17]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [18])
);
defparam \top/processor/sha_core/w[17]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [17])
);
defparam \top/processor/sha_core/w[17]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [16])
);
defparam \top/processor/sha_core/w[17]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [15])
);
defparam \top/processor/sha_core/w[17]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [14])
);
defparam \top/processor/sha_core/w[17]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [13])
);
defparam \top/processor/sha_core/w[17]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [12])
);
defparam \top/processor/sha_core/w[17]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [11])
);
defparam \top/processor/sha_core/w[17]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [10])
);
defparam \top/processor/sha_core/w[17]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [9])
);
defparam \top/processor/sha_core/w[17]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [8])
);
defparam \top/processor/sha_core/w[17]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [7])
);
defparam \top/processor/sha_core/w[17]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [6])
);
defparam \top/processor/sha_core/w[17]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [5])
);
defparam \top/processor/sha_core/w[17]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [4])
);
defparam \top/processor/sha_core/w[17]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [3])
);
defparam \top/processor/sha_core/w[17]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [2])
);
defparam \top/processor/sha_core/w[17]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [1])
);
defparam \top/processor/sha_core/w[17]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[17]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[17]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[17] [0])
);
defparam \top/processor/sha_core/w[17]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [31])
);
defparam \top/processor/sha_core/w[18]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [30])
);
defparam \top/processor/sha_core/w[18]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [29])
);
defparam \top/processor/sha_core/w[18]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [28])
);
defparam \top/processor/sha_core/w[18]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [27])
);
defparam \top/processor/sha_core/w[18]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [26])
);
defparam \top/processor/sha_core/w[18]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [25])
);
defparam \top/processor/sha_core/w[18]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [24])
);
defparam \top/processor/sha_core/w[18]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [23])
);
defparam \top/processor/sha_core/w[18]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [22])
);
defparam \top/processor/sha_core/w[18]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [21])
);
defparam \top/processor/sha_core/w[18]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [20])
);
defparam \top/processor/sha_core/w[18]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [19])
);
defparam \top/processor/sha_core/w[18]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [18])
);
defparam \top/processor/sha_core/w[18]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [17])
);
defparam \top/processor/sha_core/w[18]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [16])
);
defparam \top/processor/sha_core/w[18]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [15])
);
defparam \top/processor/sha_core/w[18]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [14])
);
defparam \top/processor/sha_core/w[18]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [13])
);
defparam \top/processor/sha_core/w[18]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [12])
);
defparam \top/processor/sha_core/w[18]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [11])
);
defparam \top/processor/sha_core/w[18]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [10])
);
defparam \top/processor/sha_core/w[18]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [9])
);
defparam \top/processor/sha_core/w[18]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [8])
);
defparam \top/processor/sha_core/w[18]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [7])
);
defparam \top/processor/sha_core/w[18]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [6])
);
defparam \top/processor/sha_core/w[18]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [5])
);
defparam \top/processor/sha_core/w[18]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [4])
);
defparam \top/processor/sha_core/w[18]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [3])
);
defparam \top/processor/sha_core/w[18]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [2])
);
defparam \top/processor/sha_core/w[18]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [1])
);
defparam \top/processor/sha_core/w[18]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[18]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[18]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[18] [0])
);
defparam \top/processor/sha_core/w[18]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [31])
);
defparam \top/processor/sha_core/w[19]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [30])
);
defparam \top/processor/sha_core/w[19]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [29])
);
defparam \top/processor/sha_core/w[19]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [28])
);
defparam \top/processor/sha_core/w[19]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [27])
);
defparam \top/processor/sha_core/w[19]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [26])
);
defparam \top/processor/sha_core/w[19]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [25])
);
defparam \top/processor/sha_core/w[19]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [24])
);
defparam \top/processor/sha_core/w[19]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [23])
);
defparam \top/processor/sha_core/w[19]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [22])
);
defparam \top/processor/sha_core/w[19]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [21])
);
defparam \top/processor/sha_core/w[19]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [20])
);
defparam \top/processor/sha_core/w[19]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [19])
);
defparam \top/processor/sha_core/w[19]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [18])
);
defparam \top/processor/sha_core/w[19]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [17])
);
defparam \top/processor/sha_core/w[19]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [16])
);
defparam \top/processor/sha_core/w[19]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [15])
);
defparam \top/processor/sha_core/w[19]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [14])
);
defparam \top/processor/sha_core/w[19]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [13])
);
defparam \top/processor/sha_core/w[19]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [12])
);
defparam \top/processor/sha_core/w[19]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [11])
);
defparam \top/processor/sha_core/w[19]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [10])
);
defparam \top/processor/sha_core/w[19]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [9])
);
defparam \top/processor/sha_core/w[19]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [8])
);
defparam \top/processor/sha_core/w[19]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [7])
);
defparam \top/processor/sha_core/w[19]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [6])
);
defparam \top/processor/sha_core/w[19]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [5])
);
defparam \top/processor/sha_core/w[19]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [4])
);
defparam \top/processor/sha_core/w[19]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [3])
);
defparam \top/processor/sha_core/w[19]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [2])
);
defparam \top/processor/sha_core/w[19]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [1])
);
defparam \top/processor/sha_core/w[19]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[19]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[19]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[19] [0])
);
defparam \top/processor/sha_core/w[19]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [31])
);
defparam \top/processor/sha_core/w[20]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [30])
);
defparam \top/processor/sha_core/w[20]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [29])
);
defparam \top/processor/sha_core/w[20]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [28])
);
defparam \top/processor/sha_core/w[20]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [27])
);
defparam \top/processor/sha_core/w[20]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [26])
);
defparam \top/processor/sha_core/w[20]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [25])
);
defparam \top/processor/sha_core/w[20]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [24])
);
defparam \top/processor/sha_core/w[20]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [23])
);
defparam \top/processor/sha_core/w[20]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [22])
);
defparam \top/processor/sha_core/w[20]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [21])
);
defparam \top/processor/sha_core/w[20]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [20])
);
defparam \top/processor/sha_core/w[20]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [19])
);
defparam \top/processor/sha_core/w[20]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [18])
);
defparam \top/processor/sha_core/w[20]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [17])
);
defparam \top/processor/sha_core/w[20]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [16])
);
defparam \top/processor/sha_core/w[20]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [15])
);
defparam \top/processor/sha_core/w[20]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [14])
);
defparam \top/processor/sha_core/w[20]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [13])
);
defparam \top/processor/sha_core/w[20]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [12])
);
defparam \top/processor/sha_core/w[20]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [11])
);
defparam \top/processor/sha_core/w[20]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [10])
);
defparam \top/processor/sha_core/w[20]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [9])
);
defparam \top/processor/sha_core/w[20]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [8])
);
defparam \top/processor/sha_core/w[20]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [7])
);
defparam \top/processor/sha_core/w[20]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [6])
);
defparam \top/processor/sha_core/w[20]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [5])
);
defparam \top/processor/sha_core/w[20]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [4])
);
defparam \top/processor/sha_core/w[20]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [3])
);
defparam \top/processor/sha_core/w[20]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [2])
);
defparam \top/processor/sha_core/w[20]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [1])
);
defparam \top/processor/sha_core/w[20]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[20]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[20]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[20] [0])
);
defparam \top/processor/sha_core/w[20]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [31])
);
defparam \top/processor/sha_core/w[21]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [30])
);
defparam \top/processor/sha_core/w[21]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [29])
);
defparam \top/processor/sha_core/w[21]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [28])
);
defparam \top/processor/sha_core/w[21]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [27])
);
defparam \top/processor/sha_core/w[21]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [26])
);
defparam \top/processor/sha_core/w[21]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [25])
);
defparam \top/processor/sha_core/w[21]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [24])
);
defparam \top/processor/sha_core/w[21]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [23])
);
defparam \top/processor/sha_core/w[21]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [22])
);
defparam \top/processor/sha_core/w[21]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [21])
);
defparam \top/processor/sha_core/w[21]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [20])
);
defparam \top/processor/sha_core/w[21]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [19])
);
defparam \top/processor/sha_core/w[21]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [18])
);
defparam \top/processor/sha_core/w[21]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [17])
);
defparam \top/processor/sha_core/w[21]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [16])
);
defparam \top/processor/sha_core/w[21]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [15])
);
defparam \top/processor/sha_core/w[21]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [14])
);
defparam \top/processor/sha_core/w[21]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [13])
);
defparam \top/processor/sha_core/w[21]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [12])
);
defparam \top/processor/sha_core/w[21]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [11])
);
defparam \top/processor/sha_core/w[21]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [10])
);
defparam \top/processor/sha_core/w[21]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [9])
);
defparam \top/processor/sha_core/w[21]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [8])
);
defparam \top/processor/sha_core/w[21]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [7])
);
defparam \top/processor/sha_core/w[21]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [6])
);
defparam \top/processor/sha_core/w[21]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [5])
);
defparam \top/processor/sha_core/w[21]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [4])
);
defparam \top/processor/sha_core/w[21]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [3])
);
defparam \top/processor/sha_core/w[21]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [2])
);
defparam \top/processor/sha_core/w[21]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [1])
);
defparam \top/processor/sha_core/w[21]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[21]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[21]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[21] [0])
);
defparam \top/processor/sha_core/w[21]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [31])
);
defparam \top/processor/sha_core/w[22]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [30])
);
defparam \top/processor/sha_core/w[22]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [29])
);
defparam \top/processor/sha_core/w[22]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [28])
);
defparam \top/processor/sha_core/w[22]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [27])
);
defparam \top/processor/sha_core/w[22]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [26])
);
defparam \top/processor/sha_core/w[22]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [25])
);
defparam \top/processor/sha_core/w[22]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [24])
);
defparam \top/processor/sha_core/w[22]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [23])
);
defparam \top/processor/sha_core/w[22]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [22])
);
defparam \top/processor/sha_core/w[22]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [21])
);
defparam \top/processor/sha_core/w[22]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [20])
);
defparam \top/processor/sha_core/w[22]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [19])
);
defparam \top/processor/sha_core/w[22]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [18])
);
defparam \top/processor/sha_core/w[22]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [17])
);
defparam \top/processor/sha_core/w[22]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [16])
);
defparam \top/processor/sha_core/w[22]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [15])
);
defparam \top/processor/sha_core/w[22]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [14])
);
defparam \top/processor/sha_core/w[22]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [13])
);
defparam \top/processor/sha_core/w[22]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [12])
);
defparam \top/processor/sha_core/w[22]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [11])
);
defparam \top/processor/sha_core/w[22]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [10])
);
defparam \top/processor/sha_core/w[22]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [9])
);
defparam \top/processor/sha_core/w[22]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [8])
);
defparam \top/processor/sha_core/w[22]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [7])
);
defparam \top/processor/sha_core/w[22]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [6])
);
defparam \top/processor/sha_core/w[22]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [5])
);
defparam \top/processor/sha_core/w[22]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [4])
);
defparam \top/processor/sha_core/w[22]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [3])
);
defparam \top/processor/sha_core/w[22]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [2])
);
defparam \top/processor/sha_core/w[22]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [1])
);
defparam \top/processor/sha_core/w[22]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[22]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[22]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[22] [0])
);
defparam \top/processor/sha_core/w[22]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [31])
);
defparam \top/processor/sha_core/w[23]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [30])
);
defparam \top/processor/sha_core/w[23]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [29])
);
defparam \top/processor/sha_core/w[23]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [28])
);
defparam \top/processor/sha_core/w[23]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [27])
);
defparam \top/processor/sha_core/w[23]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [26])
);
defparam \top/processor/sha_core/w[23]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [25])
);
defparam \top/processor/sha_core/w[23]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [24])
);
defparam \top/processor/sha_core/w[23]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [23])
);
defparam \top/processor/sha_core/w[23]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [22])
);
defparam \top/processor/sha_core/w[23]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [21])
);
defparam \top/processor/sha_core/w[23]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [20])
);
defparam \top/processor/sha_core/w[23]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [19])
);
defparam \top/processor/sha_core/w[23]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [18])
);
defparam \top/processor/sha_core/w[23]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [17])
);
defparam \top/processor/sha_core/w[23]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [16])
);
defparam \top/processor/sha_core/w[23]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [15])
);
defparam \top/processor/sha_core/w[23]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [14])
);
defparam \top/processor/sha_core/w[23]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [13])
);
defparam \top/processor/sha_core/w[23]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [12])
);
defparam \top/processor/sha_core/w[23]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [11])
);
defparam \top/processor/sha_core/w[23]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [10])
);
defparam \top/processor/sha_core/w[23]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [9])
);
defparam \top/processor/sha_core/w[23]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [8])
);
defparam \top/processor/sha_core/w[23]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [7])
);
defparam \top/processor/sha_core/w[23]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [6])
);
defparam \top/processor/sha_core/w[23]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [5])
);
defparam \top/processor/sha_core/w[23]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [4])
);
defparam \top/processor/sha_core/w[23]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [3])
);
defparam \top/processor/sha_core/w[23]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [2])
);
defparam \top/processor/sha_core/w[23]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [1])
);
defparam \top/processor/sha_core/w[23]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[23]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[23]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[23] [0])
);
defparam \top/processor/sha_core/w[23]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [31])
);
defparam \top/processor/sha_core/w[24]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [30])
);
defparam \top/processor/sha_core/w[24]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [29])
);
defparam \top/processor/sha_core/w[24]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [28])
);
defparam \top/processor/sha_core/w[24]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [27])
);
defparam \top/processor/sha_core/w[24]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [26])
);
defparam \top/processor/sha_core/w[24]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [25])
);
defparam \top/processor/sha_core/w[24]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [24])
);
defparam \top/processor/sha_core/w[24]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [23])
);
defparam \top/processor/sha_core/w[24]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [22])
);
defparam \top/processor/sha_core/w[24]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [21])
);
defparam \top/processor/sha_core/w[24]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [20])
);
defparam \top/processor/sha_core/w[24]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [19])
);
defparam \top/processor/sha_core/w[24]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [18])
);
defparam \top/processor/sha_core/w[24]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [17])
);
defparam \top/processor/sha_core/w[24]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [16])
);
defparam \top/processor/sha_core/w[24]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [15])
);
defparam \top/processor/sha_core/w[24]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [14])
);
defparam \top/processor/sha_core/w[24]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [13])
);
defparam \top/processor/sha_core/w[24]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [12])
);
defparam \top/processor/sha_core/w[24]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [11])
);
defparam \top/processor/sha_core/w[24]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [10])
);
defparam \top/processor/sha_core/w[24]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [9])
);
defparam \top/processor/sha_core/w[24]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [8])
);
defparam \top/processor/sha_core/w[24]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [7])
);
defparam \top/processor/sha_core/w[24]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [6])
);
defparam \top/processor/sha_core/w[24]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [5])
);
defparam \top/processor/sha_core/w[24]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [4])
);
defparam \top/processor/sha_core/w[24]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [3])
);
defparam \top/processor/sha_core/w[24]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [2])
);
defparam \top/processor/sha_core/w[24]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [1])
);
defparam \top/processor/sha_core/w[24]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[24]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[24]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[24] [0])
);
defparam \top/processor/sha_core/w[24]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [31])
);
defparam \top/processor/sha_core/w[25]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [30])
);
defparam \top/processor/sha_core/w[25]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [29])
);
defparam \top/processor/sha_core/w[25]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [28])
);
defparam \top/processor/sha_core/w[25]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [27])
);
defparam \top/processor/sha_core/w[25]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [26])
);
defparam \top/processor/sha_core/w[25]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [25])
);
defparam \top/processor/sha_core/w[25]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [24])
);
defparam \top/processor/sha_core/w[25]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [23])
);
defparam \top/processor/sha_core/w[25]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [22])
);
defparam \top/processor/sha_core/w[25]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [21])
);
defparam \top/processor/sha_core/w[25]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [20])
);
defparam \top/processor/sha_core/w[25]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [19])
);
defparam \top/processor/sha_core/w[25]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [18])
);
defparam \top/processor/sha_core/w[25]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [17])
);
defparam \top/processor/sha_core/w[25]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [16])
);
defparam \top/processor/sha_core/w[25]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [15])
);
defparam \top/processor/sha_core/w[25]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [14])
);
defparam \top/processor/sha_core/w[25]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [13])
);
defparam \top/processor/sha_core/w[25]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [12])
);
defparam \top/processor/sha_core/w[25]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [11])
);
defparam \top/processor/sha_core/w[25]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [10])
);
defparam \top/processor/sha_core/w[25]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [9])
);
defparam \top/processor/sha_core/w[25]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [8])
);
defparam \top/processor/sha_core/w[25]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [7])
);
defparam \top/processor/sha_core/w[25]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [6])
);
defparam \top/processor/sha_core/w[25]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [5])
);
defparam \top/processor/sha_core/w[25]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [4])
);
defparam \top/processor/sha_core/w[25]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [3])
);
defparam \top/processor/sha_core/w[25]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [2])
);
defparam \top/processor/sha_core/w[25]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [1])
);
defparam \top/processor/sha_core/w[25]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[25]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[25]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[25] [0])
);
defparam \top/processor/sha_core/w[25]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [31])
);
defparam \top/processor/sha_core/w[26]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [30])
);
defparam \top/processor/sha_core/w[26]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [29])
);
defparam \top/processor/sha_core/w[26]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [28])
);
defparam \top/processor/sha_core/w[26]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [27])
);
defparam \top/processor/sha_core/w[26]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [26])
);
defparam \top/processor/sha_core/w[26]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [25])
);
defparam \top/processor/sha_core/w[26]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [24])
);
defparam \top/processor/sha_core/w[26]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [23])
);
defparam \top/processor/sha_core/w[26]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [22])
);
defparam \top/processor/sha_core/w[26]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [21])
);
defparam \top/processor/sha_core/w[26]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [20])
);
defparam \top/processor/sha_core/w[26]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [19])
);
defparam \top/processor/sha_core/w[26]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [18])
);
defparam \top/processor/sha_core/w[26]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [17])
);
defparam \top/processor/sha_core/w[26]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [16])
);
defparam \top/processor/sha_core/w[26]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [15])
);
defparam \top/processor/sha_core/w[26]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [14])
);
defparam \top/processor/sha_core/w[26]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [13])
);
defparam \top/processor/sha_core/w[26]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [12])
);
defparam \top/processor/sha_core/w[26]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [11])
);
defparam \top/processor/sha_core/w[26]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [10])
);
defparam \top/processor/sha_core/w[26]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [9])
);
defparam \top/processor/sha_core/w[26]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [8])
);
defparam \top/processor/sha_core/w[26]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [7])
);
defparam \top/processor/sha_core/w[26]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [6])
);
defparam \top/processor/sha_core/w[26]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [5])
);
defparam \top/processor/sha_core/w[26]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [4])
);
defparam \top/processor/sha_core/w[26]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [3])
);
defparam \top/processor/sha_core/w[26]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [2])
);
defparam \top/processor/sha_core/w[26]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [1])
);
defparam \top/processor/sha_core/w[26]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[26]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[26]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[26] [0])
);
defparam \top/processor/sha_core/w[26]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [31])
);
defparam \top/processor/sha_core/w[27]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [30])
);
defparam \top/processor/sha_core/w[27]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [29])
);
defparam \top/processor/sha_core/w[27]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [28])
);
defparam \top/processor/sha_core/w[27]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [27])
);
defparam \top/processor/sha_core/w[27]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [26])
);
defparam \top/processor/sha_core/w[27]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [25])
);
defparam \top/processor/sha_core/w[27]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [24])
);
defparam \top/processor/sha_core/w[27]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [23])
);
defparam \top/processor/sha_core/w[27]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [22])
);
defparam \top/processor/sha_core/w[27]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [21])
);
defparam \top/processor/sha_core/w[27]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [20])
);
defparam \top/processor/sha_core/w[27]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [19])
);
defparam \top/processor/sha_core/w[27]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [18])
);
defparam \top/processor/sha_core/w[27]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [17])
);
defparam \top/processor/sha_core/w[27]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [16])
);
defparam \top/processor/sha_core/w[27]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [15])
);
defparam \top/processor/sha_core/w[27]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [14])
);
defparam \top/processor/sha_core/w[27]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [13])
);
defparam \top/processor/sha_core/w[27]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [12])
);
defparam \top/processor/sha_core/w[27]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [11])
);
defparam \top/processor/sha_core/w[27]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [10])
);
defparam \top/processor/sha_core/w[27]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [9])
);
defparam \top/processor/sha_core/w[27]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [8])
);
defparam \top/processor/sha_core/w[27]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [7])
);
defparam \top/processor/sha_core/w[27]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [6])
);
defparam \top/processor/sha_core/w[27]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [5])
);
defparam \top/processor/sha_core/w[27]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [4])
);
defparam \top/processor/sha_core/w[27]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [3])
);
defparam \top/processor/sha_core/w[27]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [2])
);
defparam \top/processor/sha_core/w[27]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [1])
);
defparam \top/processor/sha_core/w[27]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[27]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[27]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[27] [0])
);
defparam \top/processor/sha_core/w[27]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [31])
);
defparam \top/processor/sha_core/w[28]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [30])
);
defparam \top/processor/sha_core/w[28]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [29])
);
defparam \top/processor/sha_core/w[28]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [28])
);
defparam \top/processor/sha_core/w[28]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [27])
);
defparam \top/processor/sha_core/w[28]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [26])
);
defparam \top/processor/sha_core/w[28]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [25])
);
defparam \top/processor/sha_core/w[28]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [24])
);
defparam \top/processor/sha_core/w[28]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [23])
);
defparam \top/processor/sha_core/w[28]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [22])
);
defparam \top/processor/sha_core/w[28]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [21])
);
defparam \top/processor/sha_core/w[28]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [20])
);
defparam \top/processor/sha_core/w[28]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [19])
);
defparam \top/processor/sha_core/w[28]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [18])
);
defparam \top/processor/sha_core/w[28]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [17])
);
defparam \top/processor/sha_core/w[28]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [16])
);
defparam \top/processor/sha_core/w[28]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [15])
);
defparam \top/processor/sha_core/w[28]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [14])
);
defparam \top/processor/sha_core/w[28]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [13])
);
defparam \top/processor/sha_core/w[28]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [12])
);
defparam \top/processor/sha_core/w[28]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [11])
);
defparam \top/processor/sha_core/w[28]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [10])
);
defparam \top/processor/sha_core/w[28]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [9])
);
defparam \top/processor/sha_core/w[28]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [8])
);
defparam \top/processor/sha_core/w[28]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [7])
);
defparam \top/processor/sha_core/w[28]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [6])
);
defparam \top/processor/sha_core/w[28]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [5])
);
defparam \top/processor/sha_core/w[28]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [4])
);
defparam \top/processor/sha_core/w[28]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [3])
);
defparam \top/processor/sha_core/w[28]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [2])
);
defparam \top/processor/sha_core/w[28]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [1])
);
defparam \top/processor/sha_core/w[28]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[28]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[28]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[28] [0])
);
defparam \top/processor/sha_core/w[28]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [31])
);
defparam \top/processor/sha_core/w[29]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [30])
);
defparam \top/processor/sha_core/w[29]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [29])
);
defparam \top/processor/sha_core/w[29]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [28])
);
defparam \top/processor/sha_core/w[29]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [27])
);
defparam \top/processor/sha_core/w[29]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [26])
);
defparam \top/processor/sha_core/w[29]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [25])
);
defparam \top/processor/sha_core/w[29]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [24])
);
defparam \top/processor/sha_core/w[29]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [23])
);
defparam \top/processor/sha_core/w[29]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [22])
);
defparam \top/processor/sha_core/w[29]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [21])
);
defparam \top/processor/sha_core/w[29]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [20])
);
defparam \top/processor/sha_core/w[29]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [19])
);
defparam \top/processor/sha_core/w[29]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [18])
);
defparam \top/processor/sha_core/w[29]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [17])
);
defparam \top/processor/sha_core/w[29]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [16])
);
defparam \top/processor/sha_core/w[29]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [15])
);
defparam \top/processor/sha_core/w[29]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [14])
);
defparam \top/processor/sha_core/w[29]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [13])
);
defparam \top/processor/sha_core/w[29]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [12])
);
defparam \top/processor/sha_core/w[29]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [11])
);
defparam \top/processor/sha_core/w[29]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [10])
);
defparam \top/processor/sha_core/w[29]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [9])
);
defparam \top/processor/sha_core/w[29]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [8])
);
defparam \top/processor/sha_core/w[29]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [7])
);
defparam \top/processor/sha_core/w[29]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [6])
);
defparam \top/processor/sha_core/w[29]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [5])
);
defparam \top/processor/sha_core/w[29]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [4])
);
defparam \top/processor/sha_core/w[29]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [3])
);
defparam \top/processor/sha_core/w[29]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [2])
);
defparam \top/processor/sha_core/w[29]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [1])
);
defparam \top/processor/sha_core/w[29]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[29]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[29]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[29] [0])
);
defparam \top/processor/sha_core/w[29]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [31])
);
defparam \top/processor/sha_core/w[30]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [30])
);
defparam \top/processor/sha_core/w[30]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [29])
);
defparam \top/processor/sha_core/w[30]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [28])
);
defparam \top/processor/sha_core/w[30]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [27])
);
defparam \top/processor/sha_core/w[30]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [26])
);
defparam \top/processor/sha_core/w[30]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [25])
);
defparam \top/processor/sha_core/w[30]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [24])
);
defparam \top/processor/sha_core/w[30]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [23])
);
defparam \top/processor/sha_core/w[30]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [22])
);
defparam \top/processor/sha_core/w[30]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [21])
);
defparam \top/processor/sha_core/w[30]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [20])
);
defparam \top/processor/sha_core/w[30]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [19])
);
defparam \top/processor/sha_core/w[30]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [18])
);
defparam \top/processor/sha_core/w[30]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [17])
);
defparam \top/processor/sha_core/w[30]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [16])
);
defparam \top/processor/sha_core/w[30]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [15])
);
defparam \top/processor/sha_core/w[30]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [14])
);
defparam \top/processor/sha_core/w[30]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [13])
);
defparam \top/processor/sha_core/w[30]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [12])
);
defparam \top/processor/sha_core/w[30]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [11])
);
defparam \top/processor/sha_core/w[30]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [10])
);
defparam \top/processor/sha_core/w[30]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [9])
);
defparam \top/processor/sha_core/w[30]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [8])
);
defparam \top/processor/sha_core/w[30]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [7])
);
defparam \top/processor/sha_core/w[30]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [6])
);
defparam \top/processor/sha_core/w[30]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [5])
);
defparam \top/processor/sha_core/w[30]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [4])
);
defparam \top/processor/sha_core/w[30]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [3])
);
defparam \top/processor/sha_core/w[30]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [2])
);
defparam \top/processor/sha_core/w[30]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [1])
);
defparam \top/processor/sha_core/w[30]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[30]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[30]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[30] [0])
);
defparam \top/processor/sha_core/w[30]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [31])
);
defparam \top/processor/sha_core/w[31]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [30])
);
defparam \top/processor/sha_core/w[31]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [29])
);
defparam \top/processor/sha_core/w[31]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [28])
);
defparam \top/processor/sha_core/w[31]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [27])
);
defparam \top/processor/sha_core/w[31]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [26])
);
defparam \top/processor/sha_core/w[31]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [25])
);
defparam \top/processor/sha_core/w[31]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [24])
);
defparam \top/processor/sha_core/w[31]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [23])
);
defparam \top/processor/sha_core/w[31]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [22])
);
defparam \top/processor/sha_core/w[31]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [21])
);
defparam \top/processor/sha_core/w[31]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [20])
);
defparam \top/processor/sha_core/w[31]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [19])
);
defparam \top/processor/sha_core/w[31]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [18])
);
defparam \top/processor/sha_core/w[31]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [17])
);
defparam \top/processor/sha_core/w[31]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [16])
);
defparam \top/processor/sha_core/w[31]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [15])
);
defparam \top/processor/sha_core/w[31]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [14])
);
defparam \top/processor/sha_core/w[31]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [13])
);
defparam \top/processor/sha_core/w[31]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [12])
);
defparam \top/processor/sha_core/w[31]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [11])
);
defparam \top/processor/sha_core/w[31]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [10])
);
defparam \top/processor/sha_core/w[31]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [9])
);
defparam \top/processor/sha_core/w[31]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [8])
);
defparam \top/processor/sha_core/w[31]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [7])
);
defparam \top/processor/sha_core/w[31]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [6])
);
defparam \top/processor/sha_core/w[31]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [5])
);
defparam \top/processor/sha_core/w[31]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [4])
);
defparam \top/processor/sha_core/w[31]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [3])
);
defparam \top/processor/sha_core/w[31]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [2])
);
defparam \top/processor/sha_core/w[31]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [1])
);
defparam \top/processor/sha_core/w[31]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[31]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[31]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[31] [0])
);
defparam \top/processor/sha_core/w[31]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [31])
);
defparam \top/processor/sha_core/w[32]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [30])
);
defparam \top/processor/sha_core/w[32]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [29])
);
defparam \top/processor/sha_core/w[32]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [28])
);
defparam \top/processor/sha_core/w[32]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [27])
);
defparam \top/processor/sha_core/w[32]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [26])
);
defparam \top/processor/sha_core/w[32]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [25])
);
defparam \top/processor/sha_core/w[32]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [24])
);
defparam \top/processor/sha_core/w[32]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [23])
);
defparam \top/processor/sha_core/w[32]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [22])
);
defparam \top/processor/sha_core/w[32]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [21])
);
defparam \top/processor/sha_core/w[32]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [20])
);
defparam \top/processor/sha_core/w[32]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [19])
);
defparam \top/processor/sha_core/w[32]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [18])
);
defparam \top/processor/sha_core/w[32]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [17])
);
defparam \top/processor/sha_core/w[32]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [16])
);
defparam \top/processor/sha_core/w[32]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [15])
);
defparam \top/processor/sha_core/w[32]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [14])
);
defparam \top/processor/sha_core/w[32]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [13])
);
defparam \top/processor/sha_core/w[32]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [12])
);
defparam \top/processor/sha_core/w[32]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [11])
);
defparam \top/processor/sha_core/w[32]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [10])
);
defparam \top/processor/sha_core/w[32]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [9])
);
defparam \top/processor/sha_core/w[32]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [8])
);
defparam \top/processor/sha_core/w[32]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [7])
);
defparam \top/processor/sha_core/w[32]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [6])
);
defparam \top/processor/sha_core/w[32]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [5])
);
defparam \top/processor/sha_core/w[32]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [4])
);
defparam \top/processor/sha_core/w[32]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [3])
);
defparam \top/processor/sha_core/w[32]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [2])
);
defparam \top/processor/sha_core/w[32]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [1])
);
defparam \top/processor/sha_core/w[32]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[32]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[32]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[32] [0])
);
defparam \top/processor/sha_core/w[32]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [31])
);
defparam \top/processor/sha_core/w[33]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [30])
);
defparam \top/processor/sha_core/w[33]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [29])
);
defparam \top/processor/sha_core/w[33]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [28])
);
defparam \top/processor/sha_core/w[33]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [27])
);
defparam \top/processor/sha_core/w[33]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [26])
);
defparam \top/processor/sha_core/w[33]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [25])
);
defparam \top/processor/sha_core/w[33]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [24])
);
defparam \top/processor/sha_core/w[33]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [23])
);
defparam \top/processor/sha_core/w[33]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [22])
);
defparam \top/processor/sha_core/w[33]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [21])
);
defparam \top/processor/sha_core/w[33]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [20])
);
defparam \top/processor/sha_core/w[33]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [19])
);
defparam \top/processor/sha_core/w[33]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [18])
);
defparam \top/processor/sha_core/w[33]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [17])
);
defparam \top/processor/sha_core/w[33]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [16])
);
defparam \top/processor/sha_core/w[33]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [15])
);
defparam \top/processor/sha_core/w[33]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [14])
);
defparam \top/processor/sha_core/w[33]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [13])
);
defparam \top/processor/sha_core/w[33]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [12])
);
defparam \top/processor/sha_core/w[33]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [11])
);
defparam \top/processor/sha_core/w[33]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [10])
);
defparam \top/processor/sha_core/w[33]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [9])
);
defparam \top/processor/sha_core/w[33]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [8])
);
defparam \top/processor/sha_core/w[33]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [7])
);
defparam \top/processor/sha_core/w[33]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [6])
);
defparam \top/processor/sha_core/w[33]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [5])
);
defparam \top/processor/sha_core/w[33]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [4])
);
defparam \top/processor/sha_core/w[33]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [3])
);
defparam \top/processor/sha_core/w[33]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [2])
);
defparam \top/processor/sha_core/w[33]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [1])
);
defparam \top/processor/sha_core/w[33]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[33]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[33]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[33] [0])
);
defparam \top/processor/sha_core/w[33]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [31])
);
defparam \top/processor/sha_core/w[34]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [30])
);
defparam \top/processor/sha_core/w[34]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [29])
);
defparam \top/processor/sha_core/w[34]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [28])
);
defparam \top/processor/sha_core/w[34]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [27])
);
defparam \top/processor/sha_core/w[34]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [26])
);
defparam \top/processor/sha_core/w[34]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [25])
);
defparam \top/processor/sha_core/w[34]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [24])
);
defparam \top/processor/sha_core/w[34]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [23])
);
defparam \top/processor/sha_core/w[34]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [22])
);
defparam \top/processor/sha_core/w[34]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [21])
);
defparam \top/processor/sha_core/w[34]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [20])
);
defparam \top/processor/sha_core/w[34]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [19])
);
defparam \top/processor/sha_core/w[34]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [18])
);
defparam \top/processor/sha_core/w[34]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [17])
);
defparam \top/processor/sha_core/w[34]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [16])
);
defparam \top/processor/sha_core/w[34]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [15])
);
defparam \top/processor/sha_core/w[34]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [14])
);
defparam \top/processor/sha_core/w[34]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [13])
);
defparam \top/processor/sha_core/w[34]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [12])
);
defparam \top/processor/sha_core/w[34]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [11])
);
defparam \top/processor/sha_core/w[34]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [10])
);
defparam \top/processor/sha_core/w[34]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [9])
);
defparam \top/processor/sha_core/w[34]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [8])
);
defparam \top/processor/sha_core/w[34]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [7])
);
defparam \top/processor/sha_core/w[34]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [6])
);
defparam \top/processor/sha_core/w[34]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [5])
);
defparam \top/processor/sha_core/w[34]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [4])
);
defparam \top/processor/sha_core/w[34]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [3])
);
defparam \top/processor/sha_core/w[34]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [2])
);
defparam \top/processor/sha_core/w[34]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [1])
);
defparam \top/processor/sha_core/w[34]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[34]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[34]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[34] [0])
);
defparam \top/processor/sha_core/w[34]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [31])
);
defparam \top/processor/sha_core/w[35]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [30])
);
defparam \top/processor/sha_core/w[35]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [29])
);
defparam \top/processor/sha_core/w[35]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [28])
);
defparam \top/processor/sha_core/w[35]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [27])
);
defparam \top/processor/sha_core/w[35]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [26])
);
defparam \top/processor/sha_core/w[35]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [25])
);
defparam \top/processor/sha_core/w[35]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [24])
);
defparam \top/processor/sha_core/w[35]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [23])
);
defparam \top/processor/sha_core/w[35]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [22])
);
defparam \top/processor/sha_core/w[35]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [21])
);
defparam \top/processor/sha_core/w[35]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [20])
);
defparam \top/processor/sha_core/w[35]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [19])
);
defparam \top/processor/sha_core/w[35]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [18])
);
defparam \top/processor/sha_core/w[35]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [17])
);
defparam \top/processor/sha_core/w[35]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [16])
);
defparam \top/processor/sha_core/w[35]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [15])
);
defparam \top/processor/sha_core/w[35]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [14])
);
defparam \top/processor/sha_core/w[35]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [13])
);
defparam \top/processor/sha_core/w[35]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [12])
);
defparam \top/processor/sha_core/w[35]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [11])
);
defparam \top/processor/sha_core/w[35]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [10])
);
defparam \top/processor/sha_core/w[35]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [9])
);
defparam \top/processor/sha_core/w[35]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [8])
);
defparam \top/processor/sha_core/w[35]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [7])
);
defparam \top/processor/sha_core/w[35]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [6])
);
defparam \top/processor/sha_core/w[35]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [5])
);
defparam \top/processor/sha_core/w[35]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [4])
);
defparam \top/processor/sha_core/w[35]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [3])
);
defparam \top/processor/sha_core/w[35]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [2])
);
defparam \top/processor/sha_core/w[35]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [1])
);
defparam \top/processor/sha_core/w[35]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[35]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[35]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[35] [0])
);
defparam \top/processor/sha_core/w[35]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [31])
);
defparam \top/processor/sha_core/w[36]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [30])
);
defparam \top/processor/sha_core/w[36]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [29])
);
defparam \top/processor/sha_core/w[36]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [28])
);
defparam \top/processor/sha_core/w[36]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [27])
);
defparam \top/processor/sha_core/w[36]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [26])
);
defparam \top/processor/sha_core/w[36]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [25])
);
defparam \top/processor/sha_core/w[36]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [24])
);
defparam \top/processor/sha_core/w[36]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [23])
);
defparam \top/processor/sha_core/w[36]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [22])
);
defparam \top/processor/sha_core/w[36]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [21])
);
defparam \top/processor/sha_core/w[36]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [20])
);
defparam \top/processor/sha_core/w[36]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [19])
);
defparam \top/processor/sha_core/w[36]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [18])
);
defparam \top/processor/sha_core/w[36]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [17])
);
defparam \top/processor/sha_core/w[36]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [16])
);
defparam \top/processor/sha_core/w[36]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [15])
);
defparam \top/processor/sha_core/w[36]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [14])
);
defparam \top/processor/sha_core/w[36]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [13])
);
defparam \top/processor/sha_core/w[36]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [12])
);
defparam \top/processor/sha_core/w[36]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [11])
);
defparam \top/processor/sha_core/w[36]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [10])
);
defparam \top/processor/sha_core/w[36]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [9])
);
defparam \top/processor/sha_core/w[36]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [8])
);
defparam \top/processor/sha_core/w[36]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [7])
);
defparam \top/processor/sha_core/w[36]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [6])
);
defparam \top/processor/sha_core/w[36]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [5])
);
defparam \top/processor/sha_core/w[36]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [4])
);
defparam \top/processor/sha_core/w[36]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [3])
);
defparam \top/processor/sha_core/w[36]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [2])
);
defparam \top/processor/sha_core/w[36]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [1])
);
defparam \top/processor/sha_core/w[36]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[36]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[36]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[36] [0])
);
defparam \top/processor/sha_core/w[36]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [31])
);
defparam \top/processor/sha_core/w[37]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [30])
);
defparam \top/processor/sha_core/w[37]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [29])
);
defparam \top/processor/sha_core/w[37]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [28])
);
defparam \top/processor/sha_core/w[37]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [27])
);
defparam \top/processor/sha_core/w[37]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [26])
);
defparam \top/processor/sha_core/w[37]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [25])
);
defparam \top/processor/sha_core/w[37]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [24])
);
defparam \top/processor/sha_core/w[37]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [23])
);
defparam \top/processor/sha_core/w[37]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [22])
);
defparam \top/processor/sha_core/w[37]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [21])
);
defparam \top/processor/sha_core/w[37]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [20])
);
defparam \top/processor/sha_core/w[37]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [19])
);
defparam \top/processor/sha_core/w[37]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [18])
);
defparam \top/processor/sha_core/w[37]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [17])
);
defparam \top/processor/sha_core/w[37]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [16])
);
defparam \top/processor/sha_core/w[37]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [15])
);
defparam \top/processor/sha_core/w[37]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [14])
);
defparam \top/processor/sha_core/w[37]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [13])
);
defparam \top/processor/sha_core/w[37]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [12])
);
defparam \top/processor/sha_core/w[37]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [11])
);
defparam \top/processor/sha_core/w[37]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [10])
);
defparam \top/processor/sha_core/w[37]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [9])
);
defparam \top/processor/sha_core/w[37]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [8])
);
defparam \top/processor/sha_core/w[37]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [7])
);
defparam \top/processor/sha_core/w[37]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [6])
);
defparam \top/processor/sha_core/w[37]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [5])
);
defparam \top/processor/sha_core/w[37]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [4])
);
defparam \top/processor/sha_core/w[37]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [3])
);
defparam \top/processor/sha_core/w[37]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [2])
);
defparam \top/processor/sha_core/w[37]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [1])
);
defparam \top/processor/sha_core/w[37]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[37]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[37]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[37] [0])
);
defparam \top/processor/sha_core/w[37]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [31])
);
defparam \top/processor/sha_core/w[38]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [30])
);
defparam \top/processor/sha_core/w[38]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [29])
);
defparam \top/processor/sha_core/w[38]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [28])
);
defparam \top/processor/sha_core/w[38]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [27])
);
defparam \top/processor/sha_core/w[38]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [26])
);
defparam \top/processor/sha_core/w[38]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [25])
);
defparam \top/processor/sha_core/w[38]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [24])
);
defparam \top/processor/sha_core/w[38]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [23])
);
defparam \top/processor/sha_core/w[38]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [22])
);
defparam \top/processor/sha_core/w[38]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [21])
);
defparam \top/processor/sha_core/w[38]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [20])
);
defparam \top/processor/sha_core/w[38]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [19])
);
defparam \top/processor/sha_core/w[38]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [18])
);
defparam \top/processor/sha_core/w[38]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [17])
);
defparam \top/processor/sha_core/w[38]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [16])
);
defparam \top/processor/sha_core/w[38]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [15])
);
defparam \top/processor/sha_core/w[38]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [14])
);
defparam \top/processor/sha_core/w[38]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [13])
);
defparam \top/processor/sha_core/w[38]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [12])
);
defparam \top/processor/sha_core/w[38]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [11])
);
defparam \top/processor/sha_core/w[38]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [10])
);
defparam \top/processor/sha_core/w[38]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [9])
);
defparam \top/processor/sha_core/w[38]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [8])
);
defparam \top/processor/sha_core/w[38]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [7])
);
defparam \top/processor/sha_core/w[38]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [6])
);
defparam \top/processor/sha_core/w[38]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [5])
);
defparam \top/processor/sha_core/w[38]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [4])
);
defparam \top/processor/sha_core/w[38]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [3])
);
defparam \top/processor/sha_core/w[38]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [2])
);
defparam \top/processor/sha_core/w[38]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [1])
);
defparam \top/processor/sha_core/w[38]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[38]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[38]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[38] [0])
);
defparam \top/processor/sha_core/w[38]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [31])
);
defparam \top/processor/sha_core/w[39]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [30])
);
defparam \top/processor/sha_core/w[39]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [29])
);
defparam \top/processor/sha_core/w[39]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [28])
);
defparam \top/processor/sha_core/w[39]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [27])
);
defparam \top/processor/sha_core/w[39]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [26])
);
defparam \top/processor/sha_core/w[39]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [25])
);
defparam \top/processor/sha_core/w[39]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [24])
);
defparam \top/processor/sha_core/w[39]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [23])
);
defparam \top/processor/sha_core/w[39]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [22])
);
defparam \top/processor/sha_core/w[39]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [21])
);
defparam \top/processor/sha_core/w[39]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [20])
);
defparam \top/processor/sha_core/w[39]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [19])
);
defparam \top/processor/sha_core/w[39]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [18])
);
defparam \top/processor/sha_core/w[39]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [17])
);
defparam \top/processor/sha_core/w[39]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [16])
);
defparam \top/processor/sha_core/w[39]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [15])
);
defparam \top/processor/sha_core/w[39]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [14])
);
defparam \top/processor/sha_core/w[39]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [13])
);
defparam \top/processor/sha_core/w[39]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [12])
);
defparam \top/processor/sha_core/w[39]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [11])
);
defparam \top/processor/sha_core/w[39]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [10])
);
defparam \top/processor/sha_core/w[39]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [9])
);
defparam \top/processor/sha_core/w[39]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [8])
);
defparam \top/processor/sha_core/w[39]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [7])
);
defparam \top/processor/sha_core/w[39]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [6])
);
defparam \top/processor/sha_core/w[39]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [5])
);
defparam \top/processor/sha_core/w[39]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [4])
);
defparam \top/processor/sha_core/w[39]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [3])
);
defparam \top/processor/sha_core/w[39]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [2])
);
defparam \top/processor/sha_core/w[39]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [1])
);
defparam \top/processor/sha_core/w[39]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[39]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[39]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[39] [0])
);
defparam \top/processor/sha_core/w[39]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [31])
);
defparam \top/processor/sha_core/w[40]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [30])
);
defparam \top/processor/sha_core/w[40]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [29])
);
defparam \top/processor/sha_core/w[40]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [28])
);
defparam \top/processor/sha_core/w[40]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [27])
);
defparam \top/processor/sha_core/w[40]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [26])
);
defparam \top/processor/sha_core/w[40]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [25])
);
defparam \top/processor/sha_core/w[40]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [24])
);
defparam \top/processor/sha_core/w[40]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [23])
);
defparam \top/processor/sha_core/w[40]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [22])
);
defparam \top/processor/sha_core/w[40]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [21])
);
defparam \top/processor/sha_core/w[40]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [20])
);
defparam \top/processor/sha_core/w[40]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [19])
);
defparam \top/processor/sha_core/w[40]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [18])
);
defparam \top/processor/sha_core/w[40]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [17])
);
defparam \top/processor/sha_core/w[40]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [16])
);
defparam \top/processor/sha_core/w[40]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [15])
);
defparam \top/processor/sha_core/w[40]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [14])
);
defparam \top/processor/sha_core/w[40]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [13])
);
defparam \top/processor/sha_core/w[40]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [12])
);
defparam \top/processor/sha_core/w[40]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [11])
);
defparam \top/processor/sha_core/w[40]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [10])
);
defparam \top/processor/sha_core/w[40]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [9])
);
defparam \top/processor/sha_core/w[40]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [8])
);
defparam \top/processor/sha_core/w[40]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [7])
);
defparam \top/processor/sha_core/w[40]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [6])
);
defparam \top/processor/sha_core/w[40]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [5])
);
defparam \top/processor/sha_core/w[40]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [4])
);
defparam \top/processor/sha_core/w[40]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [3])
);
defparam \top/processor/sha_core/w[40]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [2])
);
defparam \top/processor/sha_core/w[40]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [1])
);
defparam \top/processor/sha_core/w[40]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[40]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[40]_31_11 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[40] [0])
);
defparam \top/processor/sha_core/w[40]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [31])
);
defparam \top/processor/sha_core/w[41]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [30])
);
defparam \top/processor/sha_core/w[41]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [29])
);
defparam \top/processor/sha_core/w[41]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [28])
);
defparam \top/processor/sha_core/w[41]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [27])
);
defparam \top/processor/sha_core/w[41]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [26])
);
defparam \top/processor/sha_core/w[41]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [25])
);
defparam \top/processor/sha_core/w[41]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [24])
);
defparam \top/processor/sha_core/w[41]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [23])
);
defparam \top/processor/sha_core/w[41]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [22])
);
defparam \top/processor/sha_core/w[41]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [21])
);
defparam \top/processor/sha_core/w[41]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [20])
);
defparam \top/processor/sha_core/w[41]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [19])
);
defparam \top/processor/sha_core/w[41]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [18])
);
defparam \top/processor/sha_core/w[41]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [17])
);
defparam \top/processor/sha_core/w[41]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [16])
);
defparam \top/processor/sha_core/w[41]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [15])
);
defparam \top/processor/sha_core/w[41]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [14])
);
defparam \top/processor/sha_core/w[41]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [13])
);
defparam \top/processor/sha_core/w[41]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [12])
);
defparam \top/processor/sha_core/w[41]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [11])
);
defparam \top/processor/sha_core/w[41]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [10])
);
defparam \top/processor/sha_core/w[41]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [9])
);
defparam \top/processor/sha_core/w[41]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [8])
);
defparam \top/processor/sha_core/w[41]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [7])
);
defparam \top/processor/sha_core/w[41]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [6])
);
defparam \top/processor/sha_core/w[41]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [5])
);
defparam \top/processor/sha_core/w[41]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [4])
);
defparam \top/processor/sha_core/w[41]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [3])
);
defparam \top/processor/sha_core/w[41]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [2])
);
defparam \top/processor/sha_core/w[41]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [1])
);
defparam \top/processor/sha_core/w[41]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[41]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[41]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[41] [0])
);
defparam \top/processor/sha_core/w[41]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [31])
);
defparam \top/processor/sha_core/w[42]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [30])
);
defparam \top/processor/sha_core/w[42]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [29])
);
defparam \top/processor/sha_core/w[42]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [28])
);
defparam \top/processor/sha_core/w[42]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [27])
);
defparam \top/processor/sha_core/w[42]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [26])
);
defparam \top/processor/sha_core/w[42]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [25])
);
defparam \top/processor/sha_core/w[42]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [24])
);
defparam \top/processor/sha_core/w[42]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [23])
);
defparam \top/processor/sha_core/w[42]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [22])
);
defparam \top/processor/sha_core/w[42]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [21])
);
defparam \top/processor/sha_core/w[42]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [20])
);
defparam \top/processor/sha_core/w[42]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [19])
);
defparam \top/processor/sha_core/w[42]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [18])
);
defparam \top/processor/sha_core/w[42]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [17])
);
defparam \top/processor/sha_core/w[42]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [16])
);
defparam \top/processor/sha_core/w[42]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [15])
);
defparam \top/processor/sha_core/w[42]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [14])
);
defparam \top/processor/sha_core/w[42]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [13])
);
defparam \top/processor/sha_core/w[42]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [12])
);
defparam \top/processor/sha_core/w[42]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [11])
);
defparam \top/processor/sha_core/w[42]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [10])
);
defparam \top/processor/sha_core/w[42]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [9])
);
defparam \top/processor/sha_core/w[42]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [8])
);
defparam \top/processor/sha_core/w[42]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [7])
);
defparam \top/processor/sha_core/w[42]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [6])
);
defparam \top/processor/sha_core/w[42]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [5])
);
defparam \top/processor/sha_core/w[42]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [4])
);
defparam \top/processor/sha_core/w[42]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [3])
);
defparam \top/processor/sha_core/w[42]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [2])
);
defparam \top/processor/sha_core/w[42]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [1])
);
defparam \top/processor/sha_core/w[42]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[42]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[42]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[42] [0])
);
defparam \top/processor/sha_core/w[42]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [31])
);
defparam \top/processor/sha_core/w[43]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [30])
);
defparam \top/processor/sha_core/w[43]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [29])
);
defparam \top/processor/sha_core/w[43]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [28])
);
defparam \top/processor/sha_core/w[43]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [27])
);
defparam \top/processor/sha_core/w[43]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [26])
);
defparam \top/processor/sha_core/w[43]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [25])
);
defparam \top/processor/sha_core/w[43]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [24])
);
defparam \top/processor/sha_core/w[43]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [23])
);
defparam \top/processor/sha_core/w[43]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [22])
);
defparam \top/processor/sha_core/w[43]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [21])
);
defparam \top/processor/sha_core/w[43]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [20])
);
defparam \top/processor/sha_core/w[43]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [19])
);
defparam \top/processor/sha_core/w[43]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [18])
);
defparam \top/processor/sha_core/w[43]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [17])
);
defparam \top/processor/sha_core/w[43]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [16])
);
defparam \top/processor/sha_core/w[43]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [15])
);
defparam \top/processor/sha_core/w[43]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [14])
);
defparam \top/processor/sha_core/w[43]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [13])
);
defparam \top/processor/sha_core/w[43]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [12])
);
defparam \top/processor/sha_core/w[43]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [11])
);
defparam \top/processor/sha_core/w[43]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [10])
);
defparam \top/processor/sha_core/w[43]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [9])
);
defparam \top/processor/sha_core/w[43]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [8])
);
defparam \top/processor/sha_core/w[43]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [7])
);
defparam \top/processor/sha_core/w[43]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [6])
);
defparam \top/processor/sha_core/w[43]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [5])
);
defparam \top/processor/sha_core/w[43]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [4])
);
defparam \top/processor/sha_core/w[43]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [3])
);
defparam \top/processor/sha_core/w[43]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [2])
);
defparam \top/processor/sha_core/w[43]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [1])
);
defparam \top/processor/sha_core/w[43]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[43]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[43]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[43] [0])
);
defparam \top/processor/sha_core/w[43]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [31])
);
defparam \top/processor/sha_core/w[44]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [30])
);
defparam \top/processor/sha_core/w[44]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [29])
);
defparam \top/processor/sha_core/w[44]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [28])
);
defparam \top/processor/sha_core/w[44]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [27])
);
defparam \top/processor/sha_core/w[44]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [26])
);
defparam \top/processor/sha_core/w[44]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [25])
);
defparam \top/processor/sha_core/w[44]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [24])
);
defparam \top/processor/sha_core/w[44]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [23])
);
defparam \top/processor/sha_core/w[44]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [22])
);
defparam \top/processor/sha_core/w[44]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [21])
);
defparam \top/processor/sha_core/w[44]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [20])
);
defparam \top/processor/sha_core/w[44]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [19])
);
defparam \top/processor/sha_core/w[44]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [18])
);
defparam \top/processor/sha_core/w[44]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [17])
);
defparam \top/processor/sha_core/w[44]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [16])
);
defparam \top/processor/sha_core/w[44]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [15])
);
defparam \top/processor/sha_core/w[44]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [14])
);
defparam \top/processor/sha_core/w[44]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [13])
);
defparam \top/processor/sha_core/w[44]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [12])
);
defparam \top/processor/sha_core/w[44]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [11])
);
defparam \top/processor/sha_core/w[44]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [10])
);
defparam \top/processor/sha_core/w[44]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [9])
);
defparam \top/processor/sha_core/w[44]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [8])
);
defparam \top/processor/sha_core/w[44]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [7])
);
defparam \top/processor/sha_core/w[44]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [6])
);
defparam \top/processor/sha_core/w[44]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [5])
);
defparam \top/processor/sha_core/w[44]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [4])
);
defparam \top/processor/sha_core/w[44]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [3])
);
defparam \top/processor/sha_core/w[44]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [2])
);
defparam \top/processor/sha_core/w[44]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [1])
);
defparam \top/processor/sha_core/w[44]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[44]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[44]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[44] [0])
);
defparam \top/processor/sha_core/w[44]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [31])
);
defparam \top/processor/sha_core/w[45]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [30])
);
defparam \top/processor/sha_core/w[45]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [29])
);
defparam \top/processor/sha_core/w[45]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [28])
);
defparam \top/processor/sha_core/w[45]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [27])
);
defparam \top/processor/sha_core/w[45]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [26])
);
defparam \top/processor/sha_core/w[45]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [25])
);
defparam \top/processor/sha_core/w[45]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [24])
);
defparam \top/processor/sha_core/w[45]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [23])
);
defparam \top/processor/sha_core/w[45]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [22])
);
defparam \top/processor/sha_core/w[45]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [21])
);
defparam \top/processor/sha_core/w[45]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [20])
);
defparam \top/processor/sha_core/w[45]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [19])
);
defparam \top/processor/sha_core/w[45]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [18])
);
defparam \top/processor/sha_core/w[45]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [17])
);
defparam \top/processor/sha_core/w[45]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [16])
);
defparam \top/processor/sha_core/w[45]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [15])
);
defparam \top/processor/sha_core/w[45]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [14])
);
defparam \top/processor/sha_core/w[45]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [13])
);
defparam \top/processor/sha_core/w[45]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [12])
);
defparam \top/processor/sha_core/w[45]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [11])
);
defparam \top/processor/sha_core/w[45]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [10])
);
defparam \top/processor/sha_core/w[45]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [9])
);
defparam \top/processor/sha_core/w[45]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [8])
);
defparam \top/processor/sha_core/w[45]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [7])
);
defparam \top/processor/sha_core/w[45]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [6])
);
defparam \top/processor/sha_core/w[45]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [5])
);
defparam \top/processor/sha_core/w[45]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [4])
);
defparam \top/processor/sha_core/w[45]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [3])
);
defparam \top/processor/sha_core/w[45]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [2])
);
defparam \top/processor/sha_core/w[45]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [1])
);
defparam \top/processor/sha_core/w[45]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[45]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[45]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[45] [0])
);
defparam \top/processor/sha_core/w[45]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [31])
);
defparam \top/processor/sha_core/w[46]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [30])
);
defparam \top/processor/sha_core/w[46]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [29])
);
defparam \top/processor/sha_core/w[46]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [28])
);
defparam \top/processor/sha_core/w[46]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [27])
);
defparam \top/processor/sha_core/w[46]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [26])
);
defparam \top/processor/sha_core/w[46]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [25])
);
defparam \top/processor/sha_core/w[46]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [24])
);
defparam \top/processor/sha_core/w[46]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [23])
);
defparam \top/processor/sha_core/w[46]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [22])
);
defparam \top/processor/sha_core/w[46]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [21])
);
defparam \top/processor/sha_core/w[46]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [20])
);
defparam \top/processor/sha_core/w[46]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [19])
);
defparam \top/processor/sha_core/w[46]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [18])
);
defparam \top/processor/sha_core/w[46]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [17])
);
defparam \top/processor/sha_core/w[46]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [16])
);
defparam \top/processor/sha_core/w[46]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [15])
);
defparam \top/processor/sha_core/w[46]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [14])
);
defparam \top/processor/sha_core/w[46]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [13])
);
defparam \top/processor/sha_core/w[46]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [12])
);
defparam \top/processor/sha_core/w[46]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [11])
);
defparam \top/processor/sha_core/w[46]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [10])
);
defparam \top/processor/sha_core/w[46]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [9])
);
defparam \top/processor/sha_core/w[46]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [8])
);
defparam \top/processor/sha_core/w[46]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [7])
);
defparam \top/processor/sha_core/w[46]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [6])
);
defparam \top/processor/sha_core/w[46]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [5])
);
defparam \top/processor/sha_core/w[46]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [4])
);
defparam \top/processor/sha_core/w[46]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [3])
);
defparam \top/processor/sha_core/w[46]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [2])
);
defparam \top/processor/sha_core/w[46]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [1])
);
defparam \top/processor/sha_core/w[46]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[46]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[46]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[46] [0])
);
defparam \top/processor/sha_core/w[46]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [31])
);
defparam \top/processor/sha_core/w[47]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [30])
);
defparam \top/processor/sha_core/w[47]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [29])
);
defparam \top/processor/sha_core/w[47]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [28])
);
defparam \top/processor/sha_core/w[47]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [27])
);
defparam \top/processor/sha_core/w[47]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [26])
);
defparam \top/processor/sha_core/w[47]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [25])
);
defparam \top/processor/sha_core/w[47]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [24])
);
defparam \top/processor/sha_core/w[47]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [23])
);
defparam \top/processor/sha_core/w[47]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [22])
);
defparam \top/processor/sha_core/w[47]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [21])
);
defparam \top/processor/sha_core/w[47]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [20])
);
defparam \top/processor/sha_core/w[47]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [19])
);
defparam \top/processor/sha_core/w[47]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [18])
);
defparam \top/processor/sha_core/w[47]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [17])
);
defparam \top/processor/sha_core/w[47]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [16])
);
defparam \top/processor/sha_core/w[47]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [15])
);
defparam \top/processor/sha_core/w[47]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [14])
);
defparam \top/processor/sha_core/w[47]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [13])
);
defparam \top/processor/sha_core/w[47]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [12])
);
defparam \top/processor/sha_core/w[47]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [11])
);
defparam \top/processor/sha_core/w[47]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [10])
);
defparam \top/processor/sha_core/w[47]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [9])
);
defparam \top/processor/sha_core/w[47]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [8])
);
defparam \top/processor/sha_core/w[47]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [7])
);
defparam \top/processor/sha_core/w[47]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [6])
);
defparam \top/processor/sha_core/w[47]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [5])
);
defparam \top/processor/sha_core/w[47]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [4])
);
defparam \top/processor/sha_core/w[47]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [3])
);
defparam \top/processor/sha_core/w[47]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [2])
);
defparam \top/processor/sha_core/w[47]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [1])
);
defparam \top/processor/sha_core/w[47]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[47]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[47]_31_10 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[47] [0])
);
defparam \top/processor/sha_core/w[47]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [31])
);
defparam \top/processor/sha_core/w[48]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [30])
);
defparam \top/processor/sha_core/w[48]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [29])
);
defparam \top/processor/sha_core/w[48]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [28])
);
defparam \top/processor/sha_core/w[48]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [27])
);
defparam \top/processor/sha_core/w[48]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [26])
);
defparam \top/processor/sha_core/w[48]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [25])
);
defparam \top/processor/sha_core/w[48]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [24])
);
defparam \top/processor/sha_core/w[48]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [23])
);
defparam \top/processor/sha_core/w[48]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [22])
);
defparam \top/processor/sha_core/w[48]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [21])
);
defparam \top/processor/sha_core/w[48]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [20])
);
defparam \top/processor/sha_core/w[48]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [19])
);
defparam \top/processor/sha_core/w[48]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [18])
);
defparam \top/processor/sha_core/w[48]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [17])
);
defparam \top/processor/sha_core/w[48]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [16])
);
defparam \top/processor/sha_core/w[48]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [15])
);
defparam \top/processor/sha_core/w[48]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [14])
);
defparam \top/processor/sha_core/w[48]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [13])
);
defparam \top/processor/sha_core/w[48]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [12])
);
defparam \top/processor/sha_core/w[48]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [11])
);
defparam \top/processor/sha_core/w[48]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [10])
);
defparam \top/processor/sha_core/w[48]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [9])
);
defparam \top/processor/sha_core/w[48]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [8])
);
defparam \top/processor/sha_core/w[48]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [7])
);
defparam \top/processor/sha_core/w[48]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [6])
);
defparam \top/processor/sha_core/w[48]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [5])
);
defparam \top/processor/sha_core/w[48]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [4])
);
defparam \top/processor/sha_core/w[48]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [3])
);
defparam \top/processor/sha_core/w[48]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [2])
);
defparam \top/processor/sha_core/w[48]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [1])
);
defparam \top/processor/sha_core/w[48]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[48]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[48]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[48] [0])
);
defparam \top/processor/sha_core/w[48]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [31])
);
defparam \top/processor/sha_core/w[49]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [30])
);
defparam \top/processor/sha_core/w[49]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [29])
);
defparam \top/processor/sha_core/w[49]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [28])
);
defparam \top/processor/sha_core/w[49]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [27])
);
defparam \top/processor/sha_core/w[49]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [26])
);
defparam \top/processor/sha_core/w[49]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [25])
);
defparam \top/processor/sha_core/w[49]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [24])
);
defparam \top/processor/sha_core/w[49]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [23])
);
defparam \top/processor/sha_core/w[49]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [22])
);
defparam \top/processor/sha_core/w[49]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [21])
);
defparam \top/processor/sha_core/w[49]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [20])
);
defparam \top/processor/sha_core/w[49]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [19])
);
defparam \top/processor/sha_core/w[49]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [18])
);
defparam \top/processor/sha_core/w[49]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [17])
);
defparam \top/processor/sha_core/w[49]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [16])
);
defparam \top/processor/sha_core/w[49]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [15])
);
defparam \top/processor/sha_core/w[49]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [14])
);
defparam \top/processor/sha_core/w[49]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [13])
);
defparam \top/processor/sha_core/w[49]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [12])
);
defparam \top/processor/sha_core/w[49]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [11])
);
defparam \top/processor/sha_core/w[49]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [10])
);
defparam \top/processor/sha_core/w[49]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [9])
);
defparam \top/processor/sha_core/w[49]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [8])
);
defparam \top/processor/sha_core/w[49]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [7])
);
defparam \top/processor/sha_core/w[49]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [6])
);
defparam \top/processor/sha_core/w[49]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [5])
);
defparam \top/processor/sha_core/w[49]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [4])
);
defparam \top/processor/sha_core/w[49]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [3])
);
defparam \top/processor/sha_core/w[49]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [2])
);
defparam \top/processor/sha_core/w[49]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [1])
);
defparam \top/processor/sha_core/w[49]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[49]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[49]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[49] [0])
);
defparam \top/processor/sha_core/w[49]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [31])
);
defparam \top/processor/sha_core/w[50]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [30])
);
defparam \top/processor/sha_core/w[50]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [29])
);
defparam \top/processor/sha_core/w[50]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [28])
);
defparam \top/processor/sha_core/w[50]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [27])
);
defparam \top/processor/sha_core/w[50]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [26])
);
defparam \top/processor/sha_core/w[50]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [25])
);
defparam \top/processor/sha_core/w[50]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [24])
);
defparam \top/processor/sha_core/w[50]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [23])
);
defparam \top/processor/sha_core/w[50]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [22])
);
defparam \top/processor/sha_core/w[50]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [21])
);
defparam \top/processor/sha_core/w[50]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [20])
);
defparam \top/processor/sha_core/w[50]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [19])
);
defparam \top/processor/sha_core/w[50]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [18])
);
defparam \top/processor/sha_core/w[50]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [17])
);
defparam \top/processor/sha_core/w[50]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [16])
);
defparam \top/processor/sha_core/w[50]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [15])
);
defparam \top/processor/sha_core/w[50]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [14])
);
defparam \top/processor/sha_core/w[50]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [13])
);
defparam \top/processor/sha_core/w[50]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [12])
);
defparam \top/processor/sha_core/w[50]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [11])
);
defparam \top/processor/sha_core/w[50]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [10])
);
defparam \top/processor/sha_core/w[50]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [9])
);
defparam \top/processor/sha_core/w[50]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [8])
);
defparam \top/processor/sha_core/w[50]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [7])
);
defparam \top/processor/sha_core/w[50]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [6])
);
defparam \top/processor/sha_core/w[50]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [5])
);
defparam \top/processor/sha_core/w[50]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [4])
);
defparam \top/processor/sha_core/w[50]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [3])
);
defparam \top/processor/sha_core/w[50]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [2])
);
defparam \top/processor/sha_core/w[50]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [1])
);
defparam \top/processor/sha_core/w[50]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[50]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[50]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[50] [0])
);
defparam \top/processor/sha_core/w[50]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [31])
);
defparam \top/processor/sha_core/w[51]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [30])
);
defparam \top/processor/sha_core/w[51]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [29])
);
defparam \top/processor/sha_core/w[51]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [28])
);
defparam \top/processor/sha_core/w[51]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [27])
);
defparam \top/processor/sha_core/w[51]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [26])
);
defparam \top/processor/sha_core/w[51]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [25])
);
defparam \top/processor/sha_core/w[51]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [24])
);
defparam \top/processor/sha_core/w[51]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [23])
);
defparam \top/processor/sha_core/w[51]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [22])
);
defparam \top/processor/sha_core/w[51]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [21])
);
defparam \top/processor/sha_core/w[51]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [20])
);
defparam \top/processor/sha_core/w[51]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [19])
);
defparam \top/processor/sha_core/w[51]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [18])
);
defparam \top/processor/sha_core/w[51]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [17])
);
defparam \top/processor/sha_core/w[51]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [16])
);
defparam \top/processor/sha_core/w[51]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [15])
);
defparam \top/processor/sha_core/w[51]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [14])
);
defparam \top/processor/sha_core/w[51]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [13])
);
defparam \top/processor/sha_core/w[51]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [12])
);
defparam \top/processor/sha_core/w[51]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [11])
);
defparam \top/processor/sha_core/w[51]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [10])
);
defparam \top/processor/sha_core/w[51]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [9])
);
defparam \top/processor/sha_core/w[51]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [8])
);
defparam \top/processor/sha_core/w[51]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [7])
);
defparam \top/processor/sha_core/w[51]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [6])
);
defparam \top/processor/sha_core/w[51]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [5])
);
defparam \top/processor/sha_core/w[51]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [4])
);
defparam \top/processor/sha_core/w[51]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [3])
);
defparam \top/processor/sha_core/w[51]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [2])
);
defparam \top/processor/sha_core/w[51]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [1])
);
defparam \top/processor/sha_core/w[51]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[51]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[51]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[51] [0])
);
defparam \top/processor/sha_core/w[51]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [31])
);
defparam \top/processor/sha_core/w[52]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [30])
);
defparam \top/processor/sha_core/w[52]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [29])
);
defparam \top/processor/sha_core/w[52]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [28])
);
defparam \top/processor/sha_core/w[52]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [27])
);
defparam \top/processor/sha_core/w[52]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [26])
);
defparam \top/processor/sha_core/w[52]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [25])
);
defparam \top/processor/sha_core/w[52]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [24])
);
defparam \top/processor/sha_core/w[52]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [23])
);
defparam \top/processor/sha_core/w[52]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [22])
);
defparam \top/processor/sha_core/w[52]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [21])
);
defparam \top/processor/sha_core/w[52]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [20])
);
defparam \top/processor/sha_core/w[52]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [19])
);
defparam \top/processor/sha_core/w[52]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [18])
);
defparam \top/processor/sha_core/w[52]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [17])
);
defparam \top/processor/sha_core/w[52]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [16])
);
defparam \top/processor/sha_core/w[52]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [15])
);
defparam \top/processor/sha_core/w[52]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [14])
);
defparam \top/processor/sha_core/w[52]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [13])
);
defparam \top/processor/sha_core/w[52]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [12])
);
defparam \top/processor/sha_core/w[52]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [11])
);
defparam \top/processor/sha_core/w[52]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [10])
);
defparam \top/processor/sha_core/w[52]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [9])
);
defparam \top/processor/sha_core/w[52]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [8])
);
defparam \top/processor/sha_core/w[52]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [7])
);
defparam \top/processor/sha_core/w[52]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [6])
);
defparam \top/processor/sha_core/w[52]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [5])
);
defparam \top/processor/sha_core/w[52]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [4])
);
defparam \top/processor/sha_core/w[52]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [3])
);
defparam \top/processor/sha_core/w[52]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [2])
);
defparam \top/processor/sha_core/w[52]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [1])
);
defparam \top/processor/sha_core/w[52]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[52]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[52]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[52] [0])
);
defparam \top/processor/sha_core/w[52]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [31])
);
defparam \top/processor/sha_core/w[53]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [30])
);
defparam \top/processor/sha_core/w[53]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [29])
);
defparam \top/processor/sha_core/w[53]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [28])
);
defparam \top/processor/sha_core/w[53]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [27])
);
defparam \top/processor/sha_core/w[53]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [26])
);
defparam \top/processor/sha_core/w[53]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [25])
);
defparam \top/processor/sha_core/w[53]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [24])
);
defparam \top/processor/sha_core/w[53]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [23])
);
defparam \top/processor/sha_core/w[53]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [22])
);
defparam \top/processor/sha_core/w[53]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [21])
);
defparam \top/processor/sha_core/w[53]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [20])
);
defparam \top/processor/sha_core/w[53]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [19])
);
defparam \top/processor/sha_core/w[53]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [18])
);
defparam \top/processor/sha_core/w[53]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [17])
);
defparam \top/processor/sha_core/w[53]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [16])
);
defparam \top/processor/sha_core/w[53]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [15])
);
defparam \top/processor/sha_core/w[53]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [14])
);
defparam \top/processor/sha_core/w[53]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [13])
);
defparam \top/processor/sha_core/w[53]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [12])
);
defparam \top/processor/sha_core/w[53]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [11])
);
defparam \top/processor/sha_core/w[53]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [10])
);
defparam \top/processor/sha_core/w[53]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [9])
);
defparam \top/processor/sha_core/w[53]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [8])
);
defparam \top/processor/sha_core/w[53]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [7])
);
defparam \top/processor/sha_core/w[53]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [6])
);
defparam \top/processor/sha_core/w[53]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [5])
);
defparam \top/processor/sha_core/w[53]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [4])
);
defparam \top/processor/sha_core/w[53]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [3])
);
defparam \top/processor/sha_core/w[53]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [2])
);
defparam \top/processor/sha_core/w[53]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [1])
);
defparam \top/processor/sha_core/w[53]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[53]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[53]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[53] [0])
);
defparam \top/processor/sha_core/w[53]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [31])
);
defparam \top/processor/sha_core/w[54]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [30])
);
defparam \top/processor/sha_core/w[54]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [29])
);
defparam \top/processor/sha_core/w[54]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [28])
);
defparam \top/processor/sha_core/w[54]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [27])
);
defparam \top/processor/sha_core/w[54]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [26])
);
defparam \top/processor/sha_core/w[54]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [25])
);
defparam \top/processor/sha_core/w[54]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [24])
);
defparam \top/processor/sha_core/w[54]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [23])
);
defparam \top/processor/sha_core/w[54]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [22])
);
defparam \top/processor/sha_core/w[54]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [21])
);
defparam \top/processor/sha_core/w[54]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [20])
);
defparam \top/processor/sha_core/w[54]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [19])
);
defparam \top/processor/sha_core/w[54]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [18])
);
defparam \top/processor/sha_core/w[54]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [17])
);
defparam \top/processor/sha_core/w[54]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [16])
);
defparam \top/processor/sha_core/w[54]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [15])
);
defparam \top/processor/sha_core/w[54]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [14])
);
defparam \top/processor/sha_core/w[54]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [13])
);
defparam \top/processor/sha_core/w[54]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [12])
);
defparam \top/processor/sha_core/w[54]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [11])
);
defparam \top/processor/sha_core/w[54]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [10])
);
defparam \top/processor/sha_core/w[54]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [9])
);
defparam \top/processor/sha_core/w[54]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [8])
);
defparam \top/processor/sha_core/w[54]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [7])
);
defparam \top/processor/sha_core/w[54]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [6])
);
defparam \top/processor/sha_core/w[54]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [5])
);
defparam \top/processor/sha_core/w[54]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [4])
);
defparam \top/processor/sha_core/w[54]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [3])
);
defparam \top/processor/sha_core/w[54]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [2])
);
defparam \top/processor/sha_core/w[54]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [1])
);
defparam \top/processor/sha_core/w[54]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[54]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[54]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[54] [0])
);
defparam \top/processor/sha_core/w[54]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [31])
);
defparam \top/processor/sha_core/w[55]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [30])
);
defparam \top/processor/sha_core/w[55]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [29])
);
defparam \top/processor/sha_core/w[55]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [28])
);
defparam \top/processor/sha_core/w[55]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [27])
);
defparam \top/processor/sha_core/w[55]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [26])
);
defparam \top/processor/sha_core/w[55]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [25])
);
defparam \top/processor/sha_core/w[55]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [24])
);
defparam \top/processor/sha_core/w[55]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [23])
);
defparam \top/processor/sha_core/w[55]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [22])
);
defparam \top/processor/sha_core/w[55]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [21])
);
defparam \top/processor/sha_core/w[55]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [20])
);
defparam \top/processor/sha_core/w[55]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [19])
);
defparam \top/processor/sha_core/w[55]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [18])
);
defparam \top/processor/sha_core/w[55]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [17])
);
defparam \top/processor/sha_core/w[55]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [16])
);
defparam \top/processor/sha_core/w[55]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [15])
);
defparam \top/processor/sha_core/w[55]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [14])
);
defparam \top/processor/sha_core/w[55]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [13])
);
defparam \top/processor/sha_core/w[55]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [12])
);
defparam \top/processor/sha_core/w[55]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [11])
);
defparam \top/processor/sha_core/w[55]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [10])
);
defparam \top/processor/sha_core/w[55]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [9])
);
defparam \top/processor/sha_core/w[55]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [8])
);
defparam \top/processor/sha_core/w[55]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [7])
);
defparam \top/processor/sha_core/w[55]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [6])
);
defparam \top/processor/sha_core/w[55]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [5])
);
defparam \top/processor/sha_core/w[55]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [4])
);
defparam \top/processor/sha_core/w[55]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [3])
);
defparam \top/processor/sha_core/w[55]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [2])
);
defparam \top/processor/sha_core/w[55]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [1])
);
defparam \top/processor/sha_core/w[55]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[55]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[55]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[55] [0])
);
defparam \top/processor/sha_core/w[55]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [31])
);
defparam \top/processor/sha_core/w[56]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [30])
);
defparam \top/processor/sha_core/w[56]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [29])
);
defparam \top/processor/sha_core/w[56]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [28])
);
defparam \top/processor/sha_core/w[56]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [27])
);
defparam \top/processor/sha_core/w[56]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [26])
);
defparam \top/processor/sha_core/w[56]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [25])
);
defparam \top/processor/sha_core/w[56]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [24])
);
defparam \top/processor/sha_core/w[56]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [23])
);
defparam \top/processor/sha_core/w[56]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [22])
);
defparam \top/processor/sha_core/w[56]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [21])
);
defparam \top/processor/sha_core/w[56]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [20])
);
defparam \top/processor/sha_core/w[56]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [19])
);
defparam \top/processor/sha_core/w[56]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [18])
);
defparam \top/processor/sha_core/w[56]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [17])
);
defparam \top/processor/sha_core/w[56]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [16])
);
defparam \top/processor/sha_core/w[56]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [15])
);
defparam \top/processor/sha_core/w[56]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [14])
);
defparam \top/processor/sha_core/w[56]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [13])
);
defparam \top/processor/sha_core/w[56]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [12])
);
defparam \top/processor/sha_core/w[56]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [11])
);
defparam \top/processor/sha_core/w[56]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [10])
);
defparam \top/processor/sha_core/w[56]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [9])
);
defparam \top/processor/sha_core/w[56]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [8])
);
defparam \top/processor/sha_core/w[56]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [7])
);
defparam \top/processor/sha_core/w[56]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [6])
);
defparam \top/processor/sha_core/w[56]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [5])
);
defparam \top/processor/sha_core/w[56]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [4])
);
defparam \top/processor/sha_core/w[56]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [3])
);
defparam \top/processor/sha_core/w[56]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [2])
);
defparam \top/processor/sha_core/w[56]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [1])
);
defparam \top/processor/sha_core/w[56]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[56]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[56]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[56] [0])
);
defparam \top/processor/sha_core/w[56]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [31])
);
defparam \top/processor/sha_core/w[57]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [30])
);
defparam \top/processor/sha_core/w[57]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [29])
);
defparam \top/processor/sha_core/w[57]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [28])
);
defparam \top/processor/sha_core/w[57]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [27])
);
defparam \top/processor/sha_core/w[57]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [26])
);
defparam \top/processor/sha_core/w[57]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [25])
);
defparam \top/processor/sha_core/w[57]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [24])
);
defparam \top/processor/sha_core/w[57]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [23])
);
defparam \top/processor/sha_core/w[57]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [22])
);
defparam \top/processor/sha_core/w[57]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [21])
);
defparam \top/processor/sha_core/w[57]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [20])
);
defparam \top/processor/sha_core/w[57]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [19])
);
defparam \top/processor/sha_core/w[57]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [18])
);
defparam \top/processor/sha_core/w[57]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [17])
);
defparam \top/processor/sha_core/w[57]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [16])
);
defparam \top/processor/sha_core/w[57]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [15])
);
defparam \top/processor/sha_core/w[57]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [14])
);
defparam \top/processor/sha_core/w[57]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [13])
);
defparam \top/processor/sha_core/w[57]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [12])
);
defparam \top/processor/sha_core/w[57]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [11])
);
defparam \top/processor/sha_core/w[57]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [10])
);
defparam \top/processor/sha_core/w[57]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [9])
);
defparam \top/processor/sha_core/w[57]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [8])
);
defparam \top/processor/sha_core/w[57]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [7])
);
defparam \top/processor/sha_core/w[57]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [6])
);
defparam \top/processor/sha_core/w[57]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [5])
);
defparam \top/processor/sha_core/w[57]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [4])
);
defparam \top/processor/sha_core/w[57]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [3])
);
defparam \top/processor/sha_core/w[57]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [2])
);
defparam \top/processor/sha_core/w[57]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [1])
);
defparam \top/processor/sha_core/w[57]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[57]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[57]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[57] [0])
);
defparam \top/processor/sha_core/w[57]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [31])
);
defparam \top/processor/sha_core/w[58]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [30])
);
defparam \top/processor/sha_core/w[58]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [29])
);
defparam \top/processor/sha_core/w[58]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [28])
);
defparam \top/processor/sha_core/w[58]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [27])
);
defparam \top/processor/sha_core/w[58]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [26])
);
defparam \top/processor/sha_core/w[58]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [25])
);
defparam \top/processor/sha_core/w[58]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [24])
);
defparam \top/processor/sha_core/w[58]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [23])
);
defparam \top/processor/sha_core/w[58]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [22])
);
defparam \top/processor/sha_core/w[58]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [21])
);
defparam \top/processor/sha_core/w[58]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [20])
);
defparam \top/processor/sha_core/w[58]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [19])
);
defparam \top/processor/sha_core/w[58]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [18])
);
defparam \top/processor/sha_core/w[58]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [17])
);
defparam \top/processor/sha_core/w[58]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [16])
);
defparam \top/processor/sha_core/w[58]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [15])
);
defparam \top/processor/sha_core/w[58]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [14])
);
defparam \top/processor/sha_core/w[58]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [13])
);
defparam \top/processor/sha_core/w[58]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [12])
);
defparam \top/processor/sha_core/w[58]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [11])
);
defparam \top/processor/sha_core/w[58]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [10])
);
defparam \top/processor/sha_core/w[58]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [9])
);
defparam \top/processor/sha_core/w[58]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [8])
);
defparam \top/processor/sha_core/w[58]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [7])
);
defparam \top/processor/sha_core/w[58]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [6])
);
defparam \top/processor/sha_core/w[58]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [5])
);
defparam \top/processor/sha_core/w[58]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [4])
);
defparam \top/processor/sha_core/w[58]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [3])
);
defparam \top/processor/sha_core/w[58]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [2])
);
defparam \top/processor/sha_core/w[58]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [1])
);
defparam \top/processor/sha_core/w[58]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[58]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[58]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[58] [0])
);
defparam \top/processor/sha_core/w[58]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [31])
);
defparam \top/processor/sha_core/w[59]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [30])
);
defparam \top/processor/sha_core/w[59]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [29])
);
defparam \top/processor/sha_core/w[59]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [28])
);
defparam \top/processor/sha_core/w[59]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [27])
);
defparam \top/processor/sha_core/w[59]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [26])
);
defparam \top/processor/sha_core/w[59]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [25])
);
defparam \top/processor/sha_core/w[59]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [24])
);
defparam \top/processor/sha_core/w[59]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [23])
);
defparam \top/processor/sha_core/w[59]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [22])
);
defparam \top/processor/sha_core/w[59]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [21])
);
defparam \top/processor/sha_core/w[59]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [20])
);
defparam \top/processor/sha_core/w[59]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [19])
);
defparam \top/processor/sha_core/w[59]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [18])
);
defparam \top/processor/sha_core/w[59]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [17])
);
defparam \top/processor/sha_core/w[59]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [16])
);
defparam \top/processor/sha_core/w[59]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [15])
);
defparam \top/processor/sha_core/w[59]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [14])
);
defparam \top/processor/sha_core/w[59]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [13])
);
defparam \top/processor/sha_core/w[59]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [12])
);
defparam \top/processor/sha_core/w[59]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [11])
);
defparam \top/processor/sha_core/w[59]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [10])
);
defparam \top/processor/sha_core/w[59]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [9])
);
defparam \top/processor/sha_core/w[59]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [8])
);
defparam \top/processor/sha_core/w[59]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [7])
);
defparam \top/processor/sha_core/w[59]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [6])
);
defparam \top/processor/sha_core/w[59]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [5])
);
defparam \top/processor/sha_core/w[59]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [4])
);
defparam \top/processor/sha_core/w[59]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [3])
);
defparam \top/processor/sha_core/w[59]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [2])
);
defparam \top/processor/sha_core/w[59]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [1])
);
defparam \top/processor/sha_core/w[59]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[59]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[59]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[59] [0])
);
defparam \top/processor/sha_core/w[59]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [31])
);
defparam \top/processor/sha_core/w[60]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [30])
);
defparam \top/processor/sha_core/w[60]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [29])
);
defparam \top/processor/sha_core/w[60]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [28])
);
defparam \top/processor/sha_core/w[60]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [27])
);
defparam \top/processor/sha_core/w[60]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [26])
);
defparam \top/processor/sha_core/w[60]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [25])
);
defparam \top/processor/sha_core/w[60]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [24])
);
defparam \top/processor/sha_core/w[60]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [23])
);
defparam \top/processor/sha_core/w[60]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [22])
);
defparam \top/processor/sha_core/w[60]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [21])
);
defparam \top/processor/sha_core/w[60]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [20])
);
defparam \top/processor/sha_core/w[60]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [19])
);
defparam \top/processor/sha_core/w[60]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [18])
);
defparam \top/processor/sha_core/w[60]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [17])
);
defparam \top/processor/sha_core/w[60]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [16])
);
defparam \top/processor/sha_core/w[60]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [15])
);
defparam \top/processor/sha_core/w[60]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [14])
);
defparam \top/processor/sha_core/w[60]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [13])
);
defparam \top/processor/sha_core/w[60]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [12])
);
defparam \top/processor/sha_core/w[60]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [11])
);
defparam \top/processor/sha_core/w[60]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [10])
);
defparam \top/processor/sha_core/w[60]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [9])
);
defparam \top/processor/sha_core/w[60]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [8])
);
defparam \top/processor/sha_core/w[60]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [7])
);
defparam \top/processor/sha_core/w[60]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [6])
);
defparam \top/processor/sha_core/w[60]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [5])
);
defparam \top/processor/sha_core/w[60]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [4])
);
defparam \top/processor/sha_core/w[60]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [3])
);
defparam \top/processor/sha_core/w[60]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [2])
);
defparam \top/processor/sha_core/w[60]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [1])
);
defparam \top/processor/sha_core/w[60]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[60]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[60]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[60] [0])
);
defparam \top/processor/sha_core/w[60]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [31])
);
defparam \top/processor/sha_core/w[61]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [30])
);
defparam \top/processor/sha_core/w[61]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [29])
);
defparam \top/processor/sha_core/w[61]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [28])
);
defparam \top/processor/sha_core/w[61]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [27])
);
defparam \top/processor/sha_core/w[61]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [26])
);
defparam \top/processor/sha_core/w[61]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [25])
);
defparam \top/processor/sha_core/w[61]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [24])
);
defparam \top/processor/sha_core/w[61]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [23])
);
defparam \top/processor/sha_core/w[61]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [22])
);
defparam \top/processor/sha_core/w[61]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [21])
);
defparam \top/processor/sha_core/w[61]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [20])
);
defparam \top/processor/sha_core/w[61]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [19])
);
defparam \top/processor/sha_core/w[61]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [18])
);
defparam \top/processor/sha_core/w[61]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [17])
);
defparam \top/processor/sha_core/w[61]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [16])
);
defparam \top/processor/sha_core/w[61]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [15])
);
defparam \top/processor/sha_core/w[61]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [14])
);
defparam \top/processor/sha_core/w[61]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [13])
);
defparam \top/processor/sha_core/w[61]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [12])
);
defparam \top/processor/sha_core/w[61]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [11])
);
defparam \top/processor/sha_core/w[61]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [10])
);
defparam \top/processor/sha_core/w[61]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [9])
);
defparam \top/processor/sha_core/w[61]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [8])
);
defparam \top/processor/sha_core/w[61]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [7])
);
defparam \top/processor/sha_core/w[61]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [6])
);
defparam \top/processor/sha_core/w[61]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [5])
);
defparam \top/processor/sha_core/w[61]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [4])
);
defparam \top/processor/sha_core/w[61]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [3])
);
defparam \top/processor/sha_core/w[61]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [2])
);
defparam \top/processor/sha_core/w[61]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [1])
);
defparam \top/processor/sha_core/w[61]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[61]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[61]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[61] [0])
);
defparam \top/processor/sha_core/w[61]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [31])
);
defparam \top/processor/sha_core/w[62]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [30])
);
defparam \top/processor/sha_core/w[62]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [29])
);
defparam \top/processor/sha_core/w[62]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [28])
);
defparam \top/processor/sha_core/w[62]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [27])
);
defparam \top/processor/sha_core/w[62]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [26])
);
defparam \top/processor/sha_core/w[62]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [25])
);
defparam \top/processor/sha_core/w[62]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [24])
);
defparam \top/processor/sha_core/w[62]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [23])
);
defparam \top/processor/sha_core/w[62]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [22])
);
defparam \top/processor/sha_core/w[62]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [21])
);
defparam \top/processor/sha_core/w[62]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [20])
);
defparam \top/processor/sha_core/w[62]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [19])
);
defparam \top/processor/sha_core/w[62]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [18])
);
defparam \top/processor/sha_core/w[62]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [17])
);
defparam \top/processor/sha_core/w[62]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [16])
);
defparam \top/processor/sha_core/w[62]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [15])
);
defparam \top/processor/sha_core/w[62]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [14])
);
defparam \top/processor/sha_core/w[62]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [13])
);
defparam \top/processor/sha_core/w[62]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [12])
);
defparam \top/processor/sha_core/w[62]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [11])
);
defparam \top/processor/sha_core/w[62]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [10])
);
defparam \top/processor/sha_core/w[62]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [9])
);
defparam \top/processor/sha_core/w[62]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [8])
);
defparam \top/processor/sha_core/w[62]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [7])
);
defparam \top/processor/sha_core/w[62]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [6])
);
defparam \top/processor/sha_core/w[62]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [5])
);
defparam \top/processor/sha_core/w[62]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [4])
);
defparam \top/processor/sha_core/w[62]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [3])
);
defparam \top/processor/sha_core/w[62]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [2])
);
defparam \top/processor/sha_core/w[62]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [1])
);
defparam \top/processor/sha_core/w[62]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[62]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[62]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[62] [0])
);
defparam \top/processor/sha_core/w[62]_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_31_s0  (
	.D(\top/processor/sha_core/n8430_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [31])
);
defparam \top/processor/sha_core/w[63]_31_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_30_s0  (
	.D(\top/processor/sha_core/n8431_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [30])
);
defparam \top/processor/sha_core/w[63]_30_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_29_s0  (
	.D(\top/processor/sha_core/n8432_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [29])
);
defparam \top/processor/sha_core/w[63]_29_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_28_s0  (
	.D(\top/processor/sha_core/n8433_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [28])
);
defparam \top/processor/sha_core/w[63]_28_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_27_s0  (
	.D(\top/processor/sha_core/n8434_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [27])
);
defparam \top/processor/sha_core/w[63]_27_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_26_s0  (
	.D(\top/processor/sha_core/n8435_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [26])
);
defparam \top/processor/sha_core/w[63]_26_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_25_s0  (
	.D(\top/processor/sha_core/n8436_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [25])
);
defparam \top/processor/sha_core/w[63]_25_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_24_s0  (
	.D(\top/processor/sha_core/n8437_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [24])
);
defparam \top/processor/sha_core/w[63]_24_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_23_s0  (
	.D(\top/processor/sha_core/n8438_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [23])
);
defparam \top/processor/sha_core/w[63]_23_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_22_s0  (
	.D(\top/processor/sha_core/n8439_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [22])
);
defparam \top/processor/sha_core/w[63]_22_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_21_s0  (
	.D(\top/processor/sha_core/n8440_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [21])
);
defparam \top/processor/sha_core/w[63]_21_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_20_s0  (
	.D(\top/processor/sha_core/n8441_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [20])
);
defparam \top/processor/sha_core/w[63]_20_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_19_s0  (
	.D(\top/processor/sha_core/n8442_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [19])
);
defparam \top/processor/sha_core/w[63]_19_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_18_s0  (
	.D(\top/processor/sha_core/n8443_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [18])
);
defparam \top/processor/sha_core/w[63]_18_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_17_s0  (
	.D(\top/processor/sha_core/n8444_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [17])
);
defparam \top/processor/sha_core/w[63]_17_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_16_s0  (
	.D(\top/processor/sha_core/n8445_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [16])
);
defparam \top/processor/sha_core/w[63]_16_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_15_s0  (
	.D(\top/processor/sha_core/n8446_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [15])
);
defparam \top/processor/sha_core/w[63]_15_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_14_s0  (
	.D(\top/processor/sha_core/n8447_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [14])
);
defparam \top/processor/sha_core/w[63]_14_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_13_s0  (
	.D(\top/processor/sha_core/n8448_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [13])
);
defparam \top/processor/sha_core/w[63]_13_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_12_s0  (
	.D(\top/processor/sha_core/n8449_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [12])
);
defparam \top/processor/sha_core/w[63]_12_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_11_s0  (
	.D(\top/processor/sha_core/n8450_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [11])
);
defparam \top/processor/sha_core/w[63]_11_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_10_s0  (
	.D(\top/processor/sha_core/n8451_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [10])
);
defparam \top/processor/sha_core/w[63]_10_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_9_s0  (
	.D(\top/processor/sha_core/n8452_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [9])
);
defparam \top/processor/sha_core/w[63]_9_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_8_s0  (
	.D(\top/processor/sha_core/n8453_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [8])
);
defparam \top/processor/sha_core/w[63]_8_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_7_s0  (
	.D(\top/processor/sha_core/n8454_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [7])
);
defparam \top/processor/sha_core/w[63]_7_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_6_s0  (
	.D(\top/processor/sha_core/n8455_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [6])
);
defparam \top/processor/sha_core/w[63]_6_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_5_s0  (
	.D(\top/processor/sha_core/n8456_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [5])
);
defparam \top/processor/sha_core/w[63]_5_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_4_s0  (
	.D(\top/processor/sha_core/n8457_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [4])
);
defparam \top/processor/sha_core/w[63]_4_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_3_s0  (
	.D(\top/processor/sha_core/n8458_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [3])
);
defparam \top/processor/sha_core/w[63]_3_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_2_s0  (
	.D(\top/processor/sha_core/n8459_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [2])
);
defparam \top/processor/sha_core/w[63]_2_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_1_s0  (
	.D(\top/processor/sha_core/n8460_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [1])
);
defparam \top/processor/sha_core/w[63]_1_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/w[63]_0_s0  (
	.D(\top/processor/sha_core/n8461_3 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/w[63]_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/w[63] [0])
);
defparam \top/processor/sha_core/w[63]_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_31_s0  (
	.D(\top/processor/sha_core/n11872_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [31])
);
defparam \top/processor/sha_core/h_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_30_s0  (
	.D(\top/processor/sha_core/n11873_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [30])
);
defparam \top/processor/sha_core/h_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_29_s0  (
	.D(\top/processor/sha_core/n11874_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [29])
);
defparam \top/processor/sha_core/h_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_28_s0  (
	.D(\top/processor/sha_core/n11875_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [28])
);
defparam \top/processor/sha_core/h_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_27_s0  (
	.D(\top/processor/sha_core/n11876_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [27])
);
defparam \top/processor/sha_core/h_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_26_s0  (
	.D(\top/processor/sha_core/n11877_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [26])
);
defparam \top/processor/sha_core/h_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_25_s0  (
	.D(\top/processor/sha_core/n11878_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [25])
);
defparam \top/processor/sha_core/h_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_24_s0  (
	.D(\top/processor/sha_core/n11879_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [24])
);
defparam \top/processor/sha_core/h_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_23_s0  (
	.D(\top/processor/sha_core/n11880_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [23])
);
defparam \top/processor/sha_core/h_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_22_s0  (
	.D(\top/processor/sha_core/n11881_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [22])
);
defparam \top/processor/sha_core/h_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_21_s0  (
	.D(\top/processor/sha_core/n11882_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [21])
);
defparam \top/processor/sha_core/h_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_20_s0  (
	.D(\top/processor/sha_core/n11883_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [20])
);
defparam \top/processor/sha_core/h_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_19_s0  (
	.D(\top/processor/sha_core/n11884_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [19])
);
defparam \top/processor/sha_core/h_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_18_s0  (
	.D(\top/processor/sha_core/n11885_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [18])
);
defparam \top/processor/sha_core/h_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_17_s0  (
	.D(\top/processor/sha_core/n11886_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [17])
);
defparam \top/processor/sha_core/h_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_16_s0  (
	.D(\top/processor/sha_core/n11887_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [16])
);
defparam \top/processor/sha_core/h_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_15_s0  (
	.D(\top/processor/sha_core/n11888_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [15])
);
defparam \top/processor/sha_core/h_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_14_s0  (
	.D(\top/processor/sha_core/n11889_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [14])
);
defparam \top/processor/sha_core/h_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_13_s0  (
	.D(\top/processor/sha_core/n11890_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [13])
);
defparam \top/processor/sha_core/h_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_12_s0  (
	.D(\top/processor/sha_core/n11891_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [12])
);
defparam \top/processor/sha_core/h_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_11_s0  (
	.D(\top/processor/sha_core/n11892_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [11])
);
defparam \top/processor/sha_core/h_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_10_s0  (
	.D(\top/processor/sha_core/n11893_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [10])
);
defparam \top/processor/sha_core/h_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_9_s0  (
	.D(\top/processor/sha_core/n11894_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [9])
);
defparam \top/processor/sha_core/h_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_8_s0  (
	.D(\top/processor/sha_core/n11895_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [8])
);
defparam \top/processor/sha_core/h_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_7_s0  (
	.D(\top/processor/sha_core/n11896_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [7])
);
defparam \top/processor/sha_core/h_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_6_s0  (
	.D(\top/processor/sha_core/n11897_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [6])
);
defparam \top/processor/sha_core/h_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_5_s0  (
	.D(\top/processor/sha_core/n11898_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [5])
);
defparam \top/processor/sha_core/h_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_4_s0  (
	.D(\top/processor/sha_core/n11899_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [4])
);
defparam \top/processor/sha_core/h_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_3_s0  (
	.D(\top/processor/sha_core/n11900_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [3])
);
defparam \top/processor/sha_core/h_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_2_s0  (
	.D(\top/processor/sha_core/n11901_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [2])
);
defparam \top/processor/sha_core/h_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_1_s0  (
	.D(\top/processor/sha_core/n11902_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [1])
);
defparam \top/processor/sha_core/h_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/h_0_s0  (
	.D(\top/processor/sha_core/n11903_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/h [0])
);
defparam \top/processor/sha_core/h_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_31_s0  (
	.D(\top/processor/sha_core/n11904_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [31])
);
defparam \top/processor/sha_core/g_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_30_s0  (
	.D(\top/processor/sha_core/n11905_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [30])
);
defparam \top/processor/sha_core/g_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_29_s0  (
	.D(\top/processor/sha_core/n11906_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [29])
);
defparam \top/processor/sha_core/g_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_28_s0  (
	.D(\top/processor/sha_core/n11907_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [28])
);
defparam \top/processor/sha_core/g_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_27_s0  (
	.D(\top/processor/sha_core/n11908_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [27])
);
defparam \top/processor/sha_core/g_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_26_s0  (
	.D(\top/processor/sha_core/n11909_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [26])
);
defparam \top/processor/sha_core/g_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_25_s0  (
	.D(\top/processor/sha_core/n11910_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [25])
);
defparam \top/processor/sha_core/g_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_24_s0  (
	.D(\top/processor/sha_core/n11911_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [24])
);
defparam \top/processor/sha_core/g_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_23_s0  (
	.D(\top/processor/sha_core/n11912_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [23])
);
defparam \top/processor/sha_core/g_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_22_s0  (
	.D(\top/processor/sha_core/n11913_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [22])
);
defparam \top/processor/sha_core/g_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_21_s0  (
	.D(\top/processor/sha_core/n11914_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [21])
);
defparam \top/processor/sha_core/g_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_20_s0  (
	.D(\top/processor/sha_core/n11915_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [20])
);
defparam \top/processor/sha_core/g_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_19_s0  (
	.D(\top/processor/sha_core/n11916_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [19])
);
defparam \top/processor/sha_core/g_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_18_s0  (
	.D(\top/processor/sha_core/n11917_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [18])
);
defparam \top/processor/sha_core/g_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_17_s0  (
	.D(\top/processor/sha_core/n11918_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [17])
);
defparam \top/processor/sha_core/g_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_16_s0  (
	.D(\top/processor/sha_core/n11919_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [16])
);
defparam \top/processor/sha_core/g_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_15_s0  (
	.D(\top/processor/sha_core/n11920_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [15])
);
defparam \top/processor/sha_core/g_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_14_s0  (
	.D(\top/processor/sha_core/n11921_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [14])
);
defparam \top/processor/sha_core/g_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_13_s0  (
	.D(\top/processor/sha_core/n11922_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [13])
);
defparam \top/processor/sha_core/g_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_12_s0  (
	.D(\top/processor/sha_core/n11923_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [12])
);
defparam \top/processor/sha_core/g_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_11_s0  (
	.D(\top/processor/sha_core/n11924_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [11])
);
defparam \top/processor/sha_core/g_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_10_s0  (
	.D(\top/processor/sha_core/n11925_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [10])
);
defparam \top/processor/sha_core/g_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_9_s0  (
	.D(\top/processor/sha_core/n11926_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [9])
);
defparam \top/processor/sha_core/g_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_8_s0  (
	.D(\top/processor/sha_core/n11927_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [8])
);
defparam \top/processor/sha_core/g_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_7_s0  (
	.D(\top/processor/sha_core/n11928_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [7])
);
defparam \top/processor/sha_core/g_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_6_s0  (
	.D(\top/processor/sha_core/n11929_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [6])
);
defparam \top/processor/sha_core/g_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_5_s0  (
	.D(\top/processor/sha_core/n11930_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [5])
);
defparam \top/processor/sha_core/g_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_4_s0  (
	.D(\top/processor/sha_core/n11931_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [4])
);
defparam \top/processor/sha_core/g_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_3_s0  (
	.D(\top/processor/sha_core/n11932_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [3])
);
defparam \top/processor/sha_core/g_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_2_s0  (
	.D(\top/processor/sha_core/n11933_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [2])
);
defparam \top/processor/sha_core/g_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_1_s0  (
	.D(\top/processor/sha_core/n11934_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [1])
);
defparam \top/processor/sha_core/g_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/g_0_s0  (
	.D(\top/processor/sha_core/n11935_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/g [0])
);
defparam \top/processor/sha_core/g_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_31_s0  (
	.D(\top/processor/sha_core/n11936_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [31])
);
defparam \top/processor/sha_core/f_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_30_s0  (
	.D(\top/processor/sha_core/n11937_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [30])
);
defparam \top/processor/sha_core/f_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_29_s0  (
	.D(\top/processor/sha_core/n11938_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [29])
);
defparam \top/processor/sha_core/f_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_28_s0  (
	.D(\top/processor/sha_core/n11939_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [28])
);
defparam \top/processor/sha_core/f_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_27_s0  (
	.D(\top/processor/sha_core/n11940_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [27])
);
defparam \top/processor/sha_core/f_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_26_s0  (
	.D(\top/processor/sha_core/n11941_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [26])
);
defparam \top/processor/sha_core/f_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_25_s0  (
	.D(\top/processor/sha_core/n11942_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [25])
);
defparam \top/processor/sha_core/f_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_24_s0  (
	.D(\top/processor/sha_core/n11943_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [24])
);
defparam \top/processor/sha_core/f_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_23_s0  (
	.D(\top/processor/sha_core/n11944_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [23])
);
defparam \top/processor/sha_core/f_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_22_s0  (
	.D(\top/processor/sha_core/n11945_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [22])
);
defparam \top/processor/sha_core/f_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_21_s0  (
	.D(\top/processor/sha_core/n11946_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [21])
);
defparam \top/processor/sha_core/f_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_20_s0  (
	.D(\top/processor/sha_core/n11947_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [20])
);
defparam \top/processor/sha_core/f_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_19_s0  (
	.D(\top/processor/sha_core/n11948_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [19])
);
defparam \top/processor/sha_core/f_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_18_s0  (
	.D(\top/processor/sha_core/n11949_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [18])
);
defparam \top/processor/sha_core/f_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_17_s0  (
	.D(\top/processor/sha_core/n11950_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [17])
);
defparam \top/processor/sha_core/f_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_16_s0  (
	.D(\top/processor/sha_core/n11951_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [16])
);
defparam \top/processor/sha_core/f_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_15_s0  (
	.D(\top/processor/sha_core/n11952_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [15])
);
defparam \top/processor/sha_core/f_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_14_s0  (
	.D(\top/processor/sha_core/n11953_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [14])
);
defparam \top/processor/sha_core/f_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_13_s0  (
	.D(\top/processor/sha_core/n11954_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [13])
);
defparam \top/processor/sha_core/f_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_12_s0  (
	.D(\top/processor/sha_core/n11955_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [12])
);
defparam \top/processor/sha_core/f_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_11_s0  (
	.D(\top/processor/sha_core/n11956_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [11])
);
defparam \top/processor/sha_core/f_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_10_s0  (
	.D(\top/processor/sha_core/n11957_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [10])
);
defparam \top/processor/sha_core/f_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_9_s0  (
	.D(\top/processor/sha_core/n11958_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [9])
);
defparam \top/processor/sha_core/f_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_8_s0  (
	.D(\top/processor/sha_core/n11959_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [8])
);
defparam \top/processor/sha_core/f_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_7_s0  (
	.D(\top/processor/sha_core/n11960_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [7])
);
defparam \top/processor/sha_core/f_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_6_s0  (
	.D(\top/processor/sha_core/n11961_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [6])
);
defparam \top/processor/sha_core/f_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_5_s0  (
	.D(\top/processor/sha_core/n11962_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [5])
);
defparam \top/processor/sha_core/f_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_4_s0  (
	.D(\top/processor/sha_core/n11963_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [4])
);
defparam \top/processor/sha_core/f_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_3_s0  (
	.D(\top/processor/sha_core/n11964_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [3])
);
defparam \top/processor/sha_core/f_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_2_s0  (
	.D(\top/processor/sha_core/n11965_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [2])
);
defparam \top/processor/sha_core/f_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_1_s0  (
	.D(\top/processor/sha_core/n11966_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [1])
);
defparam \top/processor/sha_core/f_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/f_0_s0  (
	.D(\top/processor/sha_core/n11967_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/f [0])
);
defparam \top/processor/sha_core/f_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_31_s0  (
	.D(\top/processor/sha_core/n11968_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [31])
);
defparam \top/processor/sha_core/e_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_30_s0  (
	.D(\top/processor/sha_core/n11969_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [30])
);
defparam \top/processor/sha_core/e_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_29_s0  (
	.D(\top/processor/sha_core/n11970_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [29])
);
defparam \top/processor/sha_core/e_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_28_s0  (
	.D(\top/processor/sha_core/n11971_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [28])
);
defparam \top/processor/sha_core/e_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_27_s0  (
	.D(\top/processor/sha_core/n11972_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [27])
);
defparam \top/processor/sha_core/e_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_26_s0  (
	.D(\top/processor/sha_core/n11973_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [26])
);
defparam \top/processor/sha_core/e_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_25_s0  (
	.D(\top/processor/sha_core/n11974_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [25])
);
defparam \top/processor/sha_core/e_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_24_s0  (
	.D(\top/processor/sha_core/n11975_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [24])
);
defparam \top/processor/sha_core/e_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_23_s0  (
	.D(\top/processor/sha_core/n11976_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [23])
);
defparam \top/processor/sha_core/e_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_22_s0  (
	.D(\top/processor/sha_core/n11977_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [22])
);
defparam \top/processor/sha_core/e_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_21_s0  (
	.D(\top/processor/sha_core/n11978_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [21])
);
defparam \top/processor/sha_core/e_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_20_s0  (
	.D(\top/processor/sha_core/n11979_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [20])
);
defparam \top/processor/sha_core/e_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_19_s0  (
	.D(\top/processor/sha_core/n11980_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [19])
);
defparam \top/processor/sha_core/e_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_18_s0  (
	.D(\top/processor/sha_core/n11981_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [18])
);
defparam \top/processor/sha_core/e_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_17_s0  (
	.D(\top/processor/sha_core/n11982_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [17])
);
defparam \top/processor/sha_core/e_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_16_s0  (
	.D(\top/processor/sha_core/n11983_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [16])
);
defparam \top/processor/sha_core/e_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_15_s0  (
	.D(\top/processor/sha_core/n11984_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [15])
);
defparam \top/processor/sha_core/e_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_14_s0  (
	.D(\top/processor/sha_core/n11985_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [14])
);
defparam \top/processor/sha_core/e_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_13_s0  (
	.D(\top/processor/sha_core/n11986_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [13])
);
defparam \top/processor/sha_core/e_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_12_s0  (
	.D(\top/processor/sha_core/n11987_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [12])
);
defparam \top/processor/sha_core/e_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_11_s0  (
	.D(\top/processor/sha_core/n11988_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [11])
);
defparam \top/processor/sha_core/e_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_10_s0  (
	.D(\top/processor/sha_core/n11989_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [10])
);
defparam \top/processor/sha_core/e_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_9_s0  (
	.D(\top/processor/sha_core/n11990_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [9])
);
defparam \top/processor/sha_core/e_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_8_s0  (
	.D(\top/processor/sha_core/n11991_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [8])
);
defparam \top/processor/sha_core/e_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_7_s0  (
	.D(\top/processor/sha_core/n11992_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [7])
);
defparam \top/processor/sha_core/e_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_6_s0  (
	.D(\top/processor/sha_core/n11993_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [6])
);
defparam \top/processor/sha_core/e_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_5_s0  (
	.D(\top/processor/sha_core/n11994_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [5])
);
defparam \top/processor/sha_core/e_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_4_s0  (
	.D(\top/processor/sha_core/n11995_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [4])
);
defparam \top/processor/sha_core/e_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_3_s0  (
	.D(\top/processor/sha_core/n11996_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [3])
);
defparam \top/processor/sha_core/e_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_2_s0  (
	.D(\top/processor/sha_core/n11997_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [2])
);
defparam \top/processor/sha_core/e_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_1_s0  (
	.D(\top/processor/sha_core/n11998_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [1])
);
defparam \top/processor/sha_core/e_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/e_0_s0  (
	.D(\top/processor/sha_core/n11999_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/e [0])
);
defparam \top/processor/sha_core/e_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_31_s0  (
	.D(\top/processor/sha_core/n12000_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [31])
);
defparam \top/processor/sha_core/d_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_30_s0  (
	.D(\top/processor/sha_core/n12001_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [30])
);
defparam \top/processor/sha_core/d_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_29_s0  (
	.D(\top/processor/sha_core/n12002_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [29])
);
defparam \top/processor/sha_core/d_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_28_s0  (
	.D(\top/processor/sha_core/n12003_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [28])
);
defparam \top/processor/sha_core/d_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_27_s0  (
	.D(\top/processor/sha_core/n12004_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [27])
);
defparam \top/processor/sha_core/d_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_26_s0  (
	.D(\top/processor/sha_core/n12005_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [26])
);
defparam \top/processor/sha_core/d_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_25_s0  (
	.D(\top/processor/sha_core/n12006_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [25])
);
defparam \top/processor/sha_core/d_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_24_s0  (
	.D(\top/processor/sha_core/n12007_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [24])
);
defparam \top/processor/sha_core/d_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_23_s0  (
	.D(\top/processor/sha_core/n12008_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [23])
);
defparam \top/processor/sha_core/d_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_22_s0  (
	.D(\top/processor/sha_core/n12009_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [22])
);
defparam \top/processor/sha_core/d_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_21_s0  (
	.D(\top/processor/sha_core/n12010_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [21])
);
defparam \top/processor/sha_core/d_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_20_s0  (
	.D(\top/processor/sha_core/n12011_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [20])
);
defparam \top/processor/sha_core/d_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_19_s0  (
	.D(\top/processor/sha_core/n12012_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [19])
);
defparam \top/processor/sha_core/d_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_18_s0  (
	.D(\top/processor/sha_core/n12013_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [18])
);
defparam \top/processor/sha_core/d_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_17_s0  (
	.D(\top/processor/sha_core/n12014_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [17])
);
defparam \top/processor/sha_core/d_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_16_s0  (
	.D(\top/processor/sha_core/n12015_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [16])
);
defparam \top/processor/sha_core/d_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_15_s0  (
	.D(\top/processor/sha_core/n12016_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [15])
);
defparam \top/processor/sha_core/d_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_14_s0  (
	.D(\top/processor/sha_core/n12017_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [14])
);
defparam \top/processor/sha_core/d_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_13_s0  (
	.D(\top/processor/sha_core/n12018_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [13])
);
defparam \top/processor/sha_core/d_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_12_s0  (
	.D(\top/processor/sha_core/n12019_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [12])
);
defparam \top/processor/sha_core/d_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_11_s0  (
	.D(\top/processor/sha_core/n12020_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [11])
);
defparam \top/processor/sha_core/d_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_10_s0  (
	.D(\top/processor/sha_core/n12021_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [10])
);
defparam \top/processor/sha_core/d_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_9_s0  (
	.D(\top/processor/sha_core/n12022_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [9])
);
defparam \top/processor/sha_core/d_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_8_s0  (
	.D(\top/processor/sha_core/n12023_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [8])
);
defparam \top/processor/sha_core/d_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_7_s0  (
	.D(\top/processor/sha_core/n12024_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [7])
);
defparam \top/processor/sha_core/d_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_6_s0  (
	.D(\top/processor/sha_core/n12025_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [6])
);
defparam \top/processor/sha_core/d_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_5_s0  (
	.D(\top/processor/sha_core/n12026_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [5])
);
defparam \top/processor/sha_core/d_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_4_s0  (
	.D(\top/processor/sha_core/n12027_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [4])
);
defparam \top/processor/sha_core/d_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_3_s0  (
	.D(\top/processor/sha_core/n12028_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [3])
);
defparam \top/processor/sha_core/d_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_2_s0  (
	.D(\top/processor/sha_core/n12029_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [2])
);
defparam \top/processor/sha_core/d_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_1_s0  (
	.D(\top/processor/sha_core/n12030_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [1])
);
defparam \top/processor/sha_core/d_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/d_0_s0  (
	.D(\top/processor/sha_core/n12031_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/d [0])
);
defparam \top/processor/sha_core/d_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_31_s0  (
	.D(\top/processor/sha_core/n12032_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [31])
);
defparam \top/processor/sha_core/c_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_30_s0  (
	.D(\top/processor/sha_core/n12033_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [30])
);
defparam \top/processor/sha_core/c_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_29_s0  (
	.D(\top/processor/sha_core/n12034_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [29])
);
defparam \top/processor/sha_core/c_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_28_s0  (
	.D(\top/processor/sha_core/n12035_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [28])
);
defparam \top/processor/sha_core/c_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_27_s0  (
	.D(\top/processor/sha_core/n12036_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [27])
);
defparam \top/processor/sha_core/c_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_26_s0  (
	.D(\top/processor/sha_core/n12037_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [26])
);
defparam \top/processor/sha_core/c_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_25_s0  (
	.D(\top/processor/sha_core/n12038_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [25])
);
defparam \top/processor/sha_core/c_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_24_s0  (
	.D(\top/processor/sha_core/n12039_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [24])
);
defparam \top/processor/sha_core/c_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_23_s0  (
	.D(\top/processor/sha_core/n12040_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [23])
);
defparam \top/processor/sha_core/c_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_22_s0  (
	.D(\top/processor/sha_core/n12041_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [22])
);
defparam \top/processor/sha_core/c_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_21_s0  (
	.D(\top/processor/sha_core/n12042_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [21])
);
defparam \top/processor/sha_core/c_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_20_s0  (
	.D(\top/processor/sha_core/n12043_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [20])
);
defparam \top/processor/sha_core/c_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_19_s0  (
	.D(\top/processor/sha_core/n12044_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [19])
);
defparam \top/processor/sha_core/c_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_18_s0  (
	.D(\top/processor/sha_core/n12045_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [18])
);
defparam \top/processor/sha_core/c_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_17_s0  (
	.D(\top/processor/sha_core/n12046_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [17])
);
defparam \top/processor/sha_core/c_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_16_s0  (
	.D(\top/processor/sha_core/n12047_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [16])
);
defparam \top/processor/sha_core/c_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_15_s0  (
	.D(\top/processor/sha_core/n12048_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [15])
);
defparam \top/processor/sha_core/c_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_14_s0  (
	.D(\top/processor/sha_core/n12049_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [14])
);
defparam \top/processor/sha_core/c_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_13_s0  (
	.D(\top/processor/sha_core/n12050_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [13])
);
defparam \top/processor/sha_core/c_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_12_s0  (
	.D(\top/processor/sha_core/n12051_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [12])
);
defparam \top/processor/sha_core/c_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_11_s0  (
	.D(\top/processor/sha_core/n12052_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [11])
);
defparam \top/processor/sha_core/c_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_10_s0  (
	.D(\top/processor/sha_core/n12053_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [10])
);
defparam \top/processor/sha_core/c_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_9_s0  (
	.D(\top/processor/sha_core/n12054_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [9])
);
defparam \top/processor/sha_core/c_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_8_s0  (
	.D(\top/processor/sha_core/n12055_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [8])
);
defparam \top/processor/sha_core/c_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_7_s0  (
	.D(\top/processor/sha_core/n12056_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [7])
);
defparam \top/processor/sha_core/c_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_6_s0  (
	.D(\top/processor/sha_core/n12057_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [6])
);
defparam \top/processor/sha_core/c_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_5_s0  (
	.D(\top/processor/sha_core/n12058_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [5])
);
defparam \top/processor/sha_core/c_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_4_s0  (
	.D(\top/processor/sha_core/n12059_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [4])
);
defparam \top/processor/sha_core/c_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_3_s0  (
	.D(\top/processor/sha_core/n12060_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [3])
);
defparam \top/processor/sha_core/c_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_2_s0  (
	.D(\top/processor/sha_core/n12061_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [2])
);
defparam \top/processor/sha_core/c_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_1_s0  (
	.D(\top/processor/sha_core/n12062_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [1])
);
defparam \top/processor/sha_core/c_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/c_0_s0  (
	.D(\top/processor/sha_core/n12063_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/c [0])
);
defparam \top/processor/sha_core/c_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_31_s0  (
	.D(\top/processor/sha_core/n12064_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [31])
);
defparam \top/processor/sha_core/b_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_30_s0  (
	.D(\top/processor/sha_core/n12065_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [30])
);
defparam \top/processor/sha_core/b_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_29_s0  (
	.D(\top/processor/sha_core/n12066_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [29])
);
defparam \top/processor/sha_core/b_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_28_s0  (
	.D(\top/processor/sha_core/n12067_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [28])
);
defparam \top/processor/sha_core/b_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_27_s0  (
	.D(\top/processor/sha_core/n12068_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [27])
);
defparam \top/processor/sha_core/b_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_26_s0  (
	.D(\top/processor/sha_core/n12069_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [26])
);
defparam \top/processor/sha_core/b_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_25_s0  (
	.D(\top/processor/sha_core/n12070_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [25])
);
defparam \top/processor/sha_core/b_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_24_s0  (
	.D(\top/processor/sha_core/n12071_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [24])
);
defparam \top/processor/sha_core/b_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_23_s0  (
	.D(\top/processor/sha_core/n12072_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [23])
);
defparam \top/processor/sha_core/b_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_22_s0  (
	.D(\top/processor/sha_core/n12073_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [22])
);
defparam \top/processor/sha_core/b_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_21_s0  (
	.D(\top/processor/sha_core/n12074_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [21])
);
defparam \top/processor/sha_core/b_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_20_s0  (
	.D(\top/processor/sha_core/n12075_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [20])
);
defparam \top/processor/sha_core/b_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_19_s0  (
	.D(\top/processor/sha_core/n12076_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [19])
);
defparam \top/processor/sha_core/b_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_18_s0  (
	.D(\top/processor/sha_core/n12077_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [18])
);
defparam \top/processor/sha_core/b_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_17_s0  (
	.D(\top/processor/sha_core/n12078_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [17])
);
defparam \top/processor/sha_core/b_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_16_s0  (
	.D(\top/processor/sha_core/n12079_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [16])
);
defparam \top/processor/sha_core/b_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_15_s0  (
	.D(\top/processor/sha_core/n12080_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [15])
);
defparam \top/processor/sha_core/b_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_14_s0  (
	.D(\top/processor/sha_core/n12081_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [14])
);
defparam \top/processor/sha_core/b_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_13_s0  (
	.D(\top/processor/sha_core/n12082_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [13])
);
defparam \top/processor/sha_core/b_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_12_s0  (
	.D(\top/processor/sha_core/n12083_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [12])
);
defparam \top/processor/sha_core/b_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_11_s0  (
	.D(\top/processor/sha_core/n12084_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [11])
);
defparam \top/processor/sha_core/b_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_10_s0  (
	.D(\top/processor/sha_core/n12085_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [10])
);
defparam \top/processor/sha_core/b_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_9_s0  (
	.D(\top/processor/sha_core/n12086_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [9])
);
defparam \top/processor/sha_core/b_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_8_s0  (
	.D(\top/processor/sha_core/n12087_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [8])
);
defparam \top/processor/sha_core/b_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_7_s0  (
	.D(\top/processor/sha_core/n12088_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [7])
);
defparam \top/processor/sha_core/b_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_6_s0  (
	.D(\top/processor/sha_core/n12089_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [6])
);
defparam \top/processor/sha_core/b_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_5_s0  (
	.D(\top/processor/sha_core/n12090_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [5])
);
defparam \top/processor/sha_core/b_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_4_s0  (
	.D(\top/processor/sha_core/n12091_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [4])
);
defparam \top/processor/sha_core/b_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_3_s0  (
	.D(\top/processor/sha_core/n12092_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [3])
);
defparam \top/processor/sha_core/b_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_2_s0  (
	.D(\top/processor/sha_core/n12093_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [2])
);
defparam \top/processor/sha_core/b_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_1_s0  (
	.D(\top/processor/sha_core/n12094_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [1])
);
defparam \top/processor/sha_core/b_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/b_0_s0  (
	.D(\top/processor/sha_core/n12095_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/b [0])
);
defparam \top/processor/sha_core/b_0_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_31_s0  (
	.D(\top/processor/sha_core/n12096_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [31])
);
defparam \top/processor/sha_core/a_31_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_30_s0  (
	.D(\top/processor/sha_core/n12097_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [30])
);
defparam \top/processor/sha_core/a_30_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_29_s0  (
	.D(\top/processor/sha_core/n12098_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [29])
);
defparam \top/processor/sha_core/a_29_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_28_s0  (
	.D(\top/processor/sha_core/n12099_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [28])
);
defparam \top/processor/sha_core/a_28_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_27_s0  (
	.D(\top/processor/sha_core/n12100_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [27])
);
defparam \top/processor/sha_core/a_27_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_26_s0  (
	.D(\top/processor/sha_core/n12101_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [26])
);
defparam \top/processor/sha_core/a_26_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_25_s0  (
	.D(\top/processor/sha_core/n12102_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [25])
);
defparam \top/processor/sha_core/a_25_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_24_s0  (
	.D(\top/processor/sha_core/n12103_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [24])
);
defparam \top/processor/sha_core/a_24_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_23_s0  (
	.D(\top/processor/sha_core/n12104_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [23])
);
defparam \top/processor/sha_core/a_23_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_22_s0  (
	.D(\top/processor/sha_core/n12105_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [22])
);
defparam \top/processor/sha_core/a_22_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_21_s0  (
	.D(\top/processor/sha_core/n12106_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [21])
);
defparam \top/processor/sha_core/a_21_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_20_s0  (
	.D(\top/processor/sha_core/n12107_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [20])
);
defparam \top/processor/sha_core/a_20_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_19_s0  (
	.D(\top/processor/sha_core/n12108_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [19])
);
defparam \top/processor/sha_core/a_19_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_18_s0  (
	.D(\top/processor/sha_core/n12109_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [18])
);
defparam \top/processor/sha_core/a_18_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_17_s0  (
	.D(\top/processor/sha_core/n12110_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [17])
);
defparam \top/processor/sha_core/a_17_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_16_s0  (
	.D(\top/processor/sha_core/n12111_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [16])
);
defparam \top/processor/sha_core/a_16_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_15_s0  (
	.D(\top/processor/sha_core/n12112_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [15])
);
defparam \top/processor/sha_core/a_15_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_14_s0  (
	.D(\top/processor/sha_core/n12113_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [14])
);
defparam \top/processor/sha_core/a_14_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_13_s0  (
	.D(\top/processor/sha_core/n12114_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [13])
);
defparam \top/processor/sha_core/a_13_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_12_s0  (
	.D(\top/processor/sha_core/n12115_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [12])
);
defparam \top/processor/sha_core/a_12_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_11_s0  (
	.D(\top/processor/sha_core/n12116_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [11])
);
defparam \top/processor/sha_core/a_11_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_10_s0  (
	.D(\top/processor/sha_core/n12117_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [10])
);
defparam \top/processor/sha_core/a_10_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_9_s0  (
	.D(\top/processor/sha_core/n12118_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [9])
);
defparam \top/processor/sha_core/a_9_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_8_s0  (
	.D(\top/processor/sha_core/n12119_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [8])
);
defparam \top/processor/sha_core/a_8_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_7_s0  (
	.D(\top/processor/sha_core/n12120_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [7])
);
defparam \top/processor/sha_core/a_7_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_6_s0  (
	.D(\top/processor/sha_core/n12121_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [6])
);
defparam \top/processor/sha_core/a_6_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_5_s0  (
	.D(\top/processor/sha_core/n12122_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [5])
);
defparam \top/processor/sha_core/a_5_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_4_s0  (
	.D(\top/processor/sha_core/n12123_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [4])
);
defparam \top/processor/sha_core/a_4_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_3_s0  (
	.D(\top/processor/sha_core/n12124_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [3])
);
defparam \top/processor/sha_core/a_3_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_2_s0  (
	.D(\top/processor/sha_core/n12125_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [2])
);
defparam \top/processor/sha_core/a_2_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_1_s0  (
	.D(\top/processor/sha_core/n12126_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [1])
);
defparam \top/processor/sha_core/a_1_s0 .INIT=1'b0;
DFFE \top/processor/sha_core/a_0_s0  (
	.D(\top/processor/sha_core/n12127_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h_31_8 ),
	.Q(\top/processor/sha_core/a [0])
);
defparam \top/processor/sha_core/a_0_s0 .INIT=1'b0;
DFFCE \top/processor/sha_core/ready_s1  (
	.D(\top/processor/sha_core/state [1]),
	.CLK(clk),
	.CE(\top/processor/sha_core/n11869_11 ),
	.CLEAR(rst),
	.Q(\top/processor/core_ready )
);
defparam \top/processor/sha_core/ready_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_6_s1  (
	.D(\top/processor/sha_core/n12128_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [6])
);
defparam \top/processor/sha_core/t_6_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_5_s1  (
	.D(\top/processor/sha_core/n12129_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [5])
);
defparam \top/processor/sha_core/t_5_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_4_s1  (
	.D(\top/processor/sha_core/n12130_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [4])
);
defparam \top/processor/sha_core/t_4_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_3_s1  (
	.D(\top/processor/sha_core/n12131_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [3])
);
defparam \top/processor/sha_core/t_3_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_2_s1  (
	.D(\top/processor/sha_core/n12132_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [2])
);
defparam \top/processor/sha_core/t_2_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_1_s1  (
	.D(\top/processor/sha_core/n12133_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [1])
);
defparam \top/processor/sha_core/t_1_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/t_0_s1  (
	.D(\top/processor/sha_core/n12134_11 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/t_6_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/t [0])
);
defparam \top/processor/sha_core/t_0_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_31_s1  (
	.D(\top/processor/sha_core/n12135_10 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [31])
);
defparam \top/processor/sha_core/h0_31_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_29_s1  (
	.D(\top/processor/sha_core/n12137_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [29])
);
defparam \top/processor/sha_core/h0_29_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_28_s1  (
	.D(\top/processor/sha_core/n12138_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [28])
);
defparam \top/processor/sha_core/h0_28_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_27_s1  (
	.D(\top/processor/sha_core/n12139_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [27])
);
defparam \top/processor/sha_core/h0_27_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_26_s1  (
	.D(\top/processor/sha_core/n12140_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [26])
);
defparam \top/processor/sha_core/h0_26_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_25_s1  (
	.D(\top/processor/sha_core/n12141_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [25])
);
defparam \top/processor/sha_core/h0_25_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_24_s1  (
	.D(\top/processor/sha_core/n12142_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [24])
);
defparam \top/processor/sha_core/h0_24_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_23_s1  (
	.D(\top/processor/sha_core/n12143_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [23])
);
defparam \top/processor/sha_core/h0_23_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_22_s1  (
	.D(\top/processor/sha_core/n12144_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [22])
);
defparam \top/processor/sha_core/h0_22_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_21_s1  (
	.D(\top/processor/sha_core/n12145_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [21])
);
defparam \top/processor/sha_core/h0_21_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_20_s1  (
	.D(\top/processor/sha_core/n12146_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [20])
);
defparam \top/processor/sha_core/h0_20_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_19_s1  (
	.D(\top/processor/sha_core/n12147_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [19])
);
defparam \top/processor/sha_core/h0_19_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_18_s1  (
	.D(\top/processor/sha_core/n12148_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [18])
);
defparam \top/processor/sha_core/h0_18_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_17_s1  (
	.D(\top/processor/sha_core/n12149_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [17])
);
defparam \top/processor/sha_core/h0_17_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_16_s1  (
	.D(\top/processor/sha_core/n12150_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [16])
);
defparam \top/processor/sha_core/h0_16_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_15_s1  (
	.D(\top/processor/sha_core/n12151_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [15])
);
defparam \top/processor/sha_core/h0_15_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_14_s1  (
	.D(\top/processor/sha_core/n12152_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [14])
);
defparam \top/processor/sha_core/h0_14_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_13_s1  (
	.D(\top/processor/sha_core/n12153_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [13])
);
defparam \top/processor/sha_core/h0_13_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_12_s1  (
	.D(\top/processor/sha_core/n12154_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [12])
);
defparam \top/processor/sha_core/h0_12_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_11_s1  (
	.D(\top/processor/sha_core/n12155_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [11])
);
defparam \top/processor/sha_core/h0_11_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_10_s1  (
	.D(\top/processor/sha_core/n12156_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [10])
);
defparam \top/processor/sha_core/h0_10_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_9_s1  (
	.D(\top/processor/sha_core/n12157_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [9])
);
defparam \top/processor/sha_core/h0_9_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_8_s1  (
	.D(\top/processor/sha_core/n12158_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [8])
);
defparam \top/processor/sha_core/h0_8_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_7_s1  (
	.D(\top/processor/sha_core/n12159_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [7])
);
defparam \top/processor/sha_core/h0_7_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_6_s1  (
	.D(\top/processor/sha_core/n12160_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [6])
);
defparam \top/processor/sha_core/h0_6_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_5_s1  (
	.D(\top/processor/sha_core/n12161_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [5])
);
defparam \top/processor/sha_core/h0_5_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h0_4_s1  (
	.D(\top/processor/sha_core/n12162_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [4])
);
defparam \top/processor/sha_core/h0_4_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h0_3_s1  (
	.D(\top/processor/sha_core/n12163_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h0 [3])
);
defparam \top/processor/sha_core/h0_3_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h0_2_s1  (
	.D(\top/processor/sha_core/n12164_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [2])
);
defparam \top/processor/sha_core/h0_2_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_1_s1  (
	.D(\top/processor/sha_core/n12165_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [1])
);
defparam \top/processor/sha_core/h0_1_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_0_s1  (
	.D(\top/processor/sha_core/n12166_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [0])
);
defparam \top/processor/sha_core/h0_0_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_31_s1  (
	.D(\top/processor/sha_core/n12167_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [31])
);
defparam \top/processor/sha_core/h1_31_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_30_s1  (
	.D(\top/processor/sha_core/n12168_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [30])
);
defparam \top/processor/sha_core/h1_30_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_29_s1  (
	.D(\top/processor/sha_core/n12169_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [29])
);
defparam \top/processor/sha_core/h1_29_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_28_s1  (
	.D(\top/processor/sha_core/n12170_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [28])
);
defparam \top/processor/sha_core/h1_28_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_27_s1  (
	.D(\top/processor/sha_core/n12171_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [27])
);
defparam \top/processor/sha_core/h1_27_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_26_s1  (
	.D(\top/processor/sha_core/n12172_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [26])
);
defparam \top/processor/sha_core/h1_26_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_25_s1  (
	.D(\top/processor/sha_core/n12173_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [25])
);
defparam \top/processor/sha_core/h1_25_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_24_s1  (
	.D(\top/processor/sha_core/n12174_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [24])
);
defparam \top/processor/sha_core/h1_24_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_23_s1  (
	.D(\top/processor/sha_core/n12175_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [23])
);
defparam \top/processor/sha_core/h1_23_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_22_s1  (
	.D(\top/processor/sha_core/n12176_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [22])
);
defparam \top/processor/sha_core/h1_22_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_21_s1  (
	.D(\top/processor/sha_core/n12177_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [21])
);
defparam \top/processor/sha_core/h1_21_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_20_s1  (
	.D(\top/processor/sha_core/n12178_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [20])
);
defparam \top/processor/sha_core/h1_20_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h1_19_s1  (
	.D(\top/processor/sha_core/n12179_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [19])
);
defparam \top/processor/sha_core/h1_19_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_18_s1  (
	.D(\top/processor/sha_core/n12180_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [18])
);
defparam \top/processor/sha_core/h1_18_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_17_s1  (
	.D(\top/processor/sha_core/n12181_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [17])
);
defparam \top/processor/sha_core/h1_17_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_16_s1  (
	.D(\top/processor/sha_core/n12182_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [16])
);
defparam \top/processor/sha_core/h1_16_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_15_s1  (
	.D(\top/processor/sha_core/n12183_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [15])
);
defparam \top/processor/sha_core/h1_15_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_14_s1  (
	.D(\top/processor/sha_core/n12184_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [14])
);
defparam \top/processor/sha_core/h1_14_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_13_s1  (
	.D(\top/processor/sha_core/n12185_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [13])
);
defparam \top/processor/sha_core/h1_13_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_12_s1  (
	.D(\top/processor/sha_core/n12186_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [12])
);
defparam \top/processor/sha_core/h1_12_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_11_s1  (
	.D(\top/processor/sha_core/n12187_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [11])
);
defparam \top/processor/sha_core/h1_11_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_10_s1  (
	.D(\top/processor/sha_core/n12188_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [10])
);
defparam \top/processor/sha_core/h1_10_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h1_9_s1  (
	.D(\top/processor/sha_core/n12189_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [9])
);
defparam \top/processor/sha_core/h1_9_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_8_s1  (
	.D(\top/processor/sha_core/n12190_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [8])
);
defparam \top/processor/sha_core/h1_8_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_7_s1  (
	.D(\top/processor/sha_core/n12191_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [7])
);
defparam \top/processor/sha_core/h1_7_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_6_s1  (
	.D(\top/processor/sha_core/n12192_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [6])
);
defparam \top/processor/sha_core/h1_6_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h1_5_s1  (
	.D(\top/processor/sha_core/n12193_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [5])
);
defparam \top/processor/sha_core/h1_5_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h1_4_s1  (
	.D(\top/processor/sha_core/n12194_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [4])
);
defparam \top/processor/sha_core/h1_4_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h1_3_s1  (
	.D(\top/processor/sha_core/n12195_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [3])
);
defparam \top/processor/sha_core/h1_3_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_2_s1  (
	.D(\top/processor/sha_core/n12196_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [2])
);
defparam \top/processor/sha_core/h1_2_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h1_1_s1  (
	.D(\top/processor/sha_core/n12197_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h1 [1])
);
defparam \top/processor/sha_core/h1_1_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h1_0_s1  (
	.D(\top/processor/sha_core/n12198_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h1 [0])
);
defparam \top/processor/sha_core/h1_0_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_31_s1  (
	.D(\top/processor/sha_core/n12199_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [31])
);
defparam \top/processor/sha_core/h2_31_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h2_30_s1  (
	.D(\top/processor/sha_core/n12200_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [30])
);
defparam \top/processor/sha_core/h2_30_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_29_s1  (
	.D(\top/processor/sha_core/n12201_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [29])
);
defparam \top/processor/sha_core/h2_29_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_28_s1  (
	.D(\top/processor/sha_core/n12202_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [28])
);
defparam \top/processor/sha_core/h2_28_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_27_s1  (
	.D(\top/processor/sha_core/n12203_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [27])
);
defparam \top/processor/sha_core/h2_27_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_26_s1  (
	.D(\top/processor/sha_core/n12204_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [26])
);
defparam \top/processor/sha_core/h2_26_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_25_s1  (
	.D(\top/processor/sha_core/n12205_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [25])
);
defparam \top/processor/sha_core/h2_25_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h2_24_s1  (
	.D(\top/processor/sha_core/n12206_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [24])
);
defparam \top/processor/sha_core/h2_24_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h2_23_s1  (
	.D(\top/processor/sha_core/n12207_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [23])
);
defparam \top/processor/sha_core/h2_23_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_22_s1  (
	.D(\top/processor/sha_core/n12208_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [22])
);
defparam \top/processor/sha_core/h2_22_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_21_s1  (
	.D(\top/processor/sha_core/n12209_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [21])
);
defparam \top/processor/sha_core/h2_21_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_20_s1  (
	.D(\top/processor/sha_core/n12210_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [20])
);
defparam \top/processor/sha_core/h2_20_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_19_s1  (
	.D(\top/processor/sha_core/n12211_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [19])
);
defparam \top/processor/sha_core/h2_19_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_18_s1  (
	.D(\top/processor/sha_core/n12212_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [18])
);
defparam \top/processor/sha_core/h2_18_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_17_s1  (
	.D(\top/processor/sha_core/n12213_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [17])
);
defparam \top/processor/sha_core/h2_17_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_16_s1  (
	.D(\top/processor/sha_core/n12214_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [16])
);
defparam \top/processor/sha_core/h2_16_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_15_s1  (
	.D(\top/processor/sha_core/n12215_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [15])
);
defparam \top/processor/sha_core/h2_15_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_14_s1  (
	.D(\top/processor/sha_core/n12216_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [14])
);
defparam \top/processor/sha_core/h2_14_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_13_s1  (
	.D(\top/processor/sha_core/n12217_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [13])
);
defparam \top/processor/sha_core/h2_13_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_12_s1  (
	.D(\top/processor/sha_core/n12218_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [12])
);
defparam \top/processor/sha_core/h2_12_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_11_s1  (
	.D(\top/processor/sha_core/n12219_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [11])
);
defparam \top/processor/sha_core/h2_11_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h2_10_s1  (
	.D(\top/processor/sha_core/n12220_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [10])
);
defparam \top/processor/sha_core/h2_10_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_9_s1  (
	.D(\top/processor/sha_core/n12221_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [9])
);
defparam \top/processor/sha_core/h2_9_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_8_s1  (
	.D(\top/processor/sha_core/n12222_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [8])
);
defparam \top/processor/sha_core/h2_8_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_7_s1  (
	.D(\top/processor/sha_core/n12223_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [7])
);
defparam \top/processor/sha_core/h2_7_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_6_s1  (
	.D(\top/processor/sha_core/n12224_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [6])
);
defparam \top/processor/sha_core/h2_6_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_5_s1  (
	.D(\top/processor/sha_core/n12225_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [5])
);
defparam \top/processor/sha_core/h2_5_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h2_4_s1  (
	.D(\top/processor/sha_core/n12226_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [4])
);
defparam \top/processor/sha_core/h2_4_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_3_s1  (
	.D(\top/processor/sha_core/n12227_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [3])
);
defparam \top/processor/sha_core/h2_3_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h2_2_s1  (
	.D(\top/processor/sha_core/n12228_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [2])
);
defparam \top/processor/sha_core/h2_2_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h2_1_s1  (
	.D(\top/processor/sha_core/n12229_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h2 [1])
);
defparam \top/processor/sha_core/h2_1_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h2_0_s1  (
	.D(\top/processor/sha_core/n12230_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h2 [0])
);
defparam \top/processor/sha_core/h2_0_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_31_s1  (
	.D(\top/processor/sha_core/n12231_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [31])
);
defparam \top/processor/sha_core/h3_31_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_30_s1  (
	.D(\top/processor/sha_core/n12232_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [30])
);
defparam \top/processor/sha_core/h3_30_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_29_s1  (
	.D(\top/processor/sha_core/n12233_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [29])
);
defparam \top/processor/sha_core/h3_29_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_28_s1  (
	.D(\top/processor/sha_core/n12234_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [28])
);
defparam \top/processor/sha_core/h3_28_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h3_27_s1  (
	.D(\top/processor/sha_core/n12235_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [27])
);
defparam \top/processor/sha_core/h3_27_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_26_s1  (
	.D(\top/processor/sha_core/n12236_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [26])
);
defparam \top/processor/sha_core/h3_26_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_25_s1  (
	.D(\top/processor/sha_core/n12237_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [25])
);
defparam \top/processor/sha_core/h3_25_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_24_s1  (
	.D(\top/processor/sha_core/n12238_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [24])
);
defparam \top/processor/sha_core/h3_24_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_23_s1  (
	.D(\top/processor/sha_core/n12239_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [23])
);
defparam \top/processor/sha_core/h3_23_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_22_s1  (
	.D(\top/processor/sha_core/n12240_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [22])
);
defparam \top/processor/sha_core/h3_22_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_21_s1  (
	.D(\top/processor/sha_core/n12241_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [21])
);
defparam \top/processor/sha_core/h3_21_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h3_20_s1  (
	.D(\top/processor/sha_core/n12242_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [20])
);
defparam \top/processor/sha_core/h3_20_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_19_s1  (
	.D(\top/processor/sha_core/n12243_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [19])
);
defparam \top/processor/sha_core/h3_19_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_18_s1  (
	.D(\top/processor/sha_core/n12244_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [18])
);
defparam \top/processor/sha_core/h3_18_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_17_s1  (
	.D(\top/processor/sha_core/n12245_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [17])
);
defparam \top/processor/sha_core/h3_17_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_16_s1  (
	.D(\top/processor/sha_core/n12246_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [16])
);
defparam \top/processor/sha_core/h3_16_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_15_s1  (
	.D(\top/processor/sha_core/n12247_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [15])
);
defparam \top/processor/sha_core/h3_15_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_14_s1  (
	.D(\top/processor/sha_core/n12248_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [14])
);
defparam \top/processor/sha_core/h3_14_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_13_s1  (
	.D(\top/processor/sha_core/n12249_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [13])
);
defparam \top/processor/sha_core/h3_13_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_12_s1  (
	.D(\top/processor/sha_core/n12250_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [12])
);
defparam \top/processor/sha_core/h3_12_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_11_s1  (
	.D(\top/processor/sha_core/n12251_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [11])
);
defparam \top/processor/sha_core/h3_11_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_10_s1  (
	.D(\top/processor/sha_core/n12252_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [10])
);
defparam \top/processor/sha_core/h3_10_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_9_s1  (
	.D(\top/processor/sha_core/n12253_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [9])
);
defparam \top/processor/sha_core/h3_9_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_8_s1  (
	.D(\top/processor/sha_core/n12254_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [8])
);
defparam \top/processor/sha_core/h3_8_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_7_s1  (
	.D(\top/processor/sha_core/n12255_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [7])
);
defparam \top/processor/sha_core/h3_7_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h3_6_s1  (
	.D(\top/processor/sha_core/n12256_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [6])
);
defparam \top/processor/sha_core/h3_6_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_5_s1  (
	.D(\top/processor/sha_core/n12257_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [5])
);
defparam \top/processor/sha_core/h3_5_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_4_s1  (
	.D(\top/processor/sha_core/n12258_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [4])
);
defparam \top/processor/sha_core/h3_4_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h3_3_s1  (
	.D(\top/processor/sha_core/n12259_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [3])
);
defparam \top/processor/sha_core/h3_3_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_2_s1  (
	.D(\top/processor/sha_core/n12260_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [2])
);
defparam \top/processor/sha_core/h3_2_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h3_1_s1  (
	.D(\top/processor/sha_core/n12261_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h3 [1])
);
defparam \top/processor/sha_core/h3_1_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h3_0_s1  (
	.D(\top/processor/sha_core/n12262_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h3 [0])
);
defparam \top/processor/sha_core/h3_0_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_31_s1  (
	.D(\top/processor/sha_core/n12263_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [31])
);
defparam \top/processor/sha_core/h4_31_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_30_s1  (
	.D(\top/processor/sha_core/n12264_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [30])
);
defparam \top/processor/sha_core/h4_30_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_29_s1  (
	.D(\top/processor/sha_core/n12265_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [29])
);
defparam \top/processor/sha_core/h4_29_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_28_s1  (
	.D(\top/processor/sha_core/n12266_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [28])
);
defparam \top/processor/sha_core/h4_28_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_27_s1  (
	.D(\top/processor/sha_core/n12267_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [27])
);
defparam \top/processor/sha_core/h4_27_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_26_s1  (
	.D(\top/processor/sha_core/n12268_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [26])
);
defparam \top/processor/sha_core/h4_26_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_25_s1  (
	.D(\top/processor/sha_core/n12269_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [25])
);
defparam \top/processor/sha_core/h4_25_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_24_s1  (
	.D(\top/processor/sha_core/n12270_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [24])
);
defparam \top/processor/sha_core/h4_24_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_23_s1  (
	.D(\top/processor/sha_core/n12271_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [23])
);
defparam \top/processor/sha_core/h4_23_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_22_s1  (
	.D(\top/processor/sha_core/n12272_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [22])
);
defparam \top/processor/sha_core/h4_22_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_21_s1  (
	.D(\top/processor/sha_core/n12273_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [21])
);
defparam \top/processor/sha_core/h4_21_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_20_s1  (
	.D(\top/processor/sha_core/n12274_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [20])
);
defparam \top/processor/sha_core/h4_20_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_19_s1  (
	.D(\top/processor/sha_core/n12275_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [19])
);
defparam \top/processor/sha_core/h4_19_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_18_s1  (
	.D(\top/processor/sha_core/n12276_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [18])
);
defparam \top/processor/sha_core/h4_18_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_17_s1  (
	.D(\top/processor/sha_core/n12277_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [17])
);
defparam \top/processor/sha_core/h4_17_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_16_s1  (
	.D(\top/processor/sha_core/n12278_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [16])
);
defparam \top/processor/sha_core/h4_16_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_15_s1  (
	.D(\top/processor/sha_core/n12279_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [15])
);
defparam \top/processor/sha_core/h4_15_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_14_s1  (
	.D(\top/processor/sha_core/n12280_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [14])
);
defparam \top/processor/sha_core/h4_14_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_13_s1  (
	.D(\top/processor/sha_core/n12281_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [13])
);
defparam \top/processor/sha_core/h4_13_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_12_s1  (
	.D(\top/processor/sha_core/n12282_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [12])
);
defparam \top/processor/sha_core/h4_12_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_11_s1  (
	.D(\top/processor/sha_core/n12283_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [11])
);
defparam \top/processor/sha_core/h4_11_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_10_s1  (
	.D(\top/processor/sha_core/n12284_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [10])
);
defparam \top/processor/sha_core/h4_10_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_9_s1  (
	.D(\top/processor/sha_core/n12285_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [9])
);
defparam \top/processor/sha_core/h4_9_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h4_8_s1  (
	.D(\top/processor/sha_core/n12286_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [8])
);
defparam \top/processor/sha_core/h4_8_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h4_7_s1  (
	.D(\top/processor/sha_core/n12287_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h4 [7])
);
defparam \top/processor/sha_core/h4_7_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h4_6_s1  (
	.D(\top/processor/sha_core/n12288_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [6])
);
defparam \top/processor/sha_core/h4_6_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_5_s1  (
	.D(\top/processor/sha_core/n12289_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [5])
);
defparam \top/processor/sha_core/h4_5_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_4_s1  (
	.D(\top/processor/sha_core/n12290_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [4])
);
defparam \top/processor/sha_core/h4_4_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_3_s1  (
	.D(\top/processor/sha_core/n12291_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [3])
);
defparam \top/processor/sha_core/h4_3_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_2_s1  (
	.D(\top/processor/sha_core/n12292_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [2])
);
defparam \top/processor/sha_core/h4_2_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_1_s1  (
	.D(\top/processor/sha_core/n12293_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [1])
);
defparam \top/processor/sha_core/h4_1_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h4_0_s1  (
	.D(\top/processor/sha_core/n12294_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h4 [0])
);
defparam \top/processor/sha_core/h4_0_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h5_31_s1  (
	.D(\top/processor/sha_core/n12295_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [31])
);
defparam \top/processor/sha_core/h5_31_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_30_s1  (
	.D(\top/processor/sha_core/n12296_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [30])
);
defparam \top/processor/sha_core/h5_30_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_29_s1  (
	.D(\top/processor/sha_core/n12297_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [29])
);
defparam \top/processor/sha_core/h5_29_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_28_s1  (
	.D(\top/processor/sha_core/n12298_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [28])
);
defparam \top/processor/sha_core/h5_28_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h5_27_s1  (
	.D(\top/processor/sha_core/n12299_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [27])
);
defparam \top/processor/sha_core/h5_27_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_26_s1  (
	.D(\top/processor/sha_core/n12300_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [26])
);
defparam \top/processor/sha_core/h5_26_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_25_s1  (
	.D(\top/processor/sha_core/n12301_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [25])
);
defparam \top/processor/sha_core/h5_25_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h5_24_s1  (
	.D(\top/processor/sha_core/n12302_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [24])
);
defparam \top/processor/sha_core/h5_24_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_23_s1  (
	.D(\top/processor/sha_core/n12303_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [23])
);
defparam \top/processor/sha_core/h5_23_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_22_s1  (
	.D(\top/processor/sha_core/n12304_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [22])
);
defparam \top/processor/sha_core/h5_22_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_21_s1  (
	.D(\top/processor/sha_core/n12305_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [21])
);
defparam \top/processor/sha_core/h5_21_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_20_s1  (
	.D(\top/processor/sha_core/n12306_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [20])
);
defparam \top/processor/sha_core/h5_20_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_19_s1  (
	.D(\top/processor/sha_core/n12307_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [19])
);
defparam \top/processor/sha_core/h5_19_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_18_s1  (
	.D(\top/processor/sha_core/n12308_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [18])
);
defparam \top/processor/sha_core/h5_18_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_17_s1  (
	.D(\top/processor/sha_core/n12309_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [17])
);
defparam \top/processor/sha_core/h5_17_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_16_s1  (
	.D(\top/processor/sha_core/n12310_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [16])
);
defparam \top/processor/sha_core/h5_16_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_15_s1  (
	.D(\top/processor/sha_core/n12311_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [15])
);
defparam \top/processor/sha_core/h5_15_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_14_s1  (
	.D(\top/processor/sha_core/n12312_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [14])
);
defparam \top/processor/sha_core/h5_14_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h5_13_s1  (
	.D(\top/processor/sha_core/n12313_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [13])
);
defparam \top/processor/sha_core/h5_13_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_12_s1  (
	.D(\top/processor/sha_core/n12314_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [12])
);
defparam \top/processor/sha_core/h5_12_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_11_s1  (
	.D(\top/processor/sha_core/n12315_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [11])
);
defparam \top/processor/sha_core/h5_11_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_10_s1  (
	.D(\top/processor/sha_core/n12316_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [10])
);
defparam \top/processor/sha_core/h5_10_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_9_s1  (
	.D(\top/processor/sha_core/n12317_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [9])
);
defparam \top/processor/sha_core/h5_9_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_8_s1  (
	.D(\top/processor/sha_core/n12318_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [8])
);
defparam \top/processor/sha_core/h5_8_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_7_s1  (
	.D(\top/processor/sha_core/n12319_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [7])
);
defparam \top/processor/sha_core/h5_7_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_6_s1  (
	.D(\top/processor/sha_core/n12320_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [6])
);
defparam \top/processor/sha_core/h5_6_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_5_s1  (
	.D(\top/processor/sha_core/n12321_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [5])
);
defparam \top/processor/sha_core/h5_5_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_4_s1  (
	.D(\top/processor/sha_core/n12322_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [4])
);
defparam \top/processor/sha_core/h5_4_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h5_3_s1  (
	.D(\top/processor/sha_core/n12323_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [3])
);
defparam \top/processor/sha_core/h5_3_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h5_2_s1  (
	.D(\top/processor/sha_core/n12324_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h5 [2])
);
defparam \top/processor/sha_core/h5_2_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h5_1_s1  (
	.D(\top/processor/sha_core/n12325_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [1])
);
defparam \top/processor/sha_core/h5_1_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h5_0_s1  (
	.D(\top/processor/sha_core/n12326_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h5 [0])
);
defparam \top/processor/sha_core/h5_0_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_31_s1  (
	.D(\top/processor/sha_core/n12327_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [31])
);
defparam \top/processor/sha_core/h6_31_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_30_s1  (
	.D(\top/processor/sha_core/n12328_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [30])
);
defparam \top/processor/sha_core/h6_30_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_29_s1  (
	.D(\top/processor/sha_core/n12329_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [29])
);
defparam \top/processor/sha_core/h6_29_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_28_s1  (
	.D(\top/processor/sha_core/n12330_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [28])
);
defparam \top/processor/sha_core/h6_28_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_27_s1  (
	.D(\top/processor/sha_core/n12331_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [27])
);
defparam \top/processor/sha_core/h6_27_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_26_s1  (
	.D(\top/processor/sha_core/n12332_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [26])
);
defparam \top/processor/sha_core/h6_26_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_25_s1  (
	.D(\top/processor/sha_core/n12333_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [25])
);
defparam \top/processor/sha_core/h6_25_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_24_s1  (
	.D(\top/processor/sha_core/n12334_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [24])
);
defparam \top/processor/sha_core/h6_24_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_23_s1  (
	.D(\top/processor/sha_core/n12335_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [23])
);
defparam \top/processor/sha_core/h6_23_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h6_22_s1  (
	.D(\top/processor/sha_core/n12336_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [22])
);
defparam \top/processor/sha_core/h6_22_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_21_s1  (
	.D(\top/processor/sha_core/n12337_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [21])
);
defparam \top/processor/sha_core/h6_21_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_20_s1  (
	.D(\top/processor/sha_core/n12338_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [20])
);
defparam \top/processor/sha_core/h6_20_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_19_s1  (
	.D(\top/processor/sha_core/n12339_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [19])
);
defparam \top/processor/sha_core/h6_19_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_18_s1  (
	.D(\top/processor/sha_core/n12340_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [18])
);
defparam \top/processor/sha_core/h6_18_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_17_s1  (
	.D(\top/processor/sha_core/n12341_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [17])
);
defparam \top/processor/sha_core/h6_17_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_16_s1  (
	.D(\top/processor/sha_core/n12342_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [16])
);
defparam \top/processor/sha_core/h6_16_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_15_s1  (
	.D(\top/processor/sha_core/n12343_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [15])
);
defparam \top/processor/sha_core/h6_15_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_14_s1  (
	.D(\top/processor/sha_core/n12344_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [14])
);
defparam \top/processor/sha_core/h6_14_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h6_13_s1  (
	.D(\top/processor/sha_core/n12345_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [13])
);
defparam \top/processor/sha_core/h6_13_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_12_s1  (
	.D(\top/processor/sha_core/n12346_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [12])
);
defparam \top/processor/sha_core/h6_12_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_11_s1  (
	.D(\top/processor/sha_core/n12347_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [11])
);
defparam \top/processor/sha_core/h6_11_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h6_10_s1  (
	.D(\top/processor/sha_core/n12348_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [10])
);
defparam \top/processor/sha_core/h6_10_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h6_9_s1  (
	.D(\top/processor/sha_core/n12349_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [9])
);
defparam \top/processor/sha_core/h6_9_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_8_s1  (
	.D(\top/processor/sha_core/n12350_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [8])
);
defparam \top/processor/sha_core/h6_8_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_7_s1  (
	.D(\top/processor/sha_core/n12351_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [7])
);
defparam \top/processor/sha_core/h6_7_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h6_6_s1  (
	.D(\top/processor/sha_core/n12352_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [6])
);
defparam \top/processor/sha_core/h6_6_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_5_s1  (
	.D(\top/processor/sha_core/n12353_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [5])
);
defparam \top/processor/sha_core/h6_5_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h6_4_s1  (
	.D(\top/processor/sha_core/n12354_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [4])
);
defparam \top/processor/sha_core/h6_4_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_3_s1  (
	.D(\top/processor/sha_core/n12355_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [3])
);
defparam \top/processor/sha_core/h6_3_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h6_2_s1  (
	.D(\top/processor/sha_core/n12356_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h6 [2])
);
defparam \top/processor/sha_core/h6_2_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h6_1_s1  (
	.D(\top/processor/sha_core/n12357_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [1])
);
defparam \top/processor/sha_core/h6_1_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h6_0_s1  (
	.D(\top/processor/sha_core/n12358_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h6 [0])
);
defparam \top/processor/sha_core/h6_0_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_31_s1  (
	.D(\top/processor/sha_core/n12359_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [31])
);
defparam \top/processor/sha_core/h7_31_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_30_s1  (
	.D(\top/processor/sha_core/n12360_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [30])
);
defparam \top/processor/sha_core/h7_30_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_29_s1  (
	.D(\top/processor/sha_core/n12361_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [29])
);
defparam \top/processor/sha_core/h7_29_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_28_s1  (
	.D(\top/processor/sha_core/n12362_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [28])
);
defparam \top/processor/sha_core/h7_28_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_27_s1  (
	.D(\top/processor/sha_core/n12363_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [27])
);
defparam \top/processor/sha_core/h7_27_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_26_s1  (
	.D(\top/processor/sha_core/n12364_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [26])
);
defparam \top/processor/sha_core/h7_26_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_25_s1  (
	.D(\top/processor/sha_core/n12365_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [25])
);
defparam \top/processor/sha_core/h7_25_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_24_s1  (
	.D(\top/processor/sha_core/n12366_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [24])
);
defparam \top/processor/sha_core/h7_24_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_23_s1  (
	.D(\top/processor/sha_core/n12367_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [23])
);
defparam \top/processor/sha_core/h7_23_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_22_s1  (
	.D(\top/processor/sha_core/n12368_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [22])
);
defparam \top/processor/sha_core/h7_22_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_21_s1  (
	.D(\top/processor/sha_core/n12369_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [21])
);
defparam \top/processor/sha_core/h7_21_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_20_s1  (
	.D(\top/processor/sha_core/n12370_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [20])
);
defparam \top/processor/sha_core/h7_20_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_19_s1  (
	.D(\top/processor/sha_core/n12371_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [19])
);
defparam \top/processor/sha_core/h7_19_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_18_s1  (
	.D(\top/processor/sha_core/n12372_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [18])
);
defparam \top/processor/sha_core/h7_18_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_17_s1  (
	.D(\top/processor/sha_core/n12373_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [17])
);
defparam \top/processor/sha_core/h7_17_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_16_s1  (
	.D(\top/processor/sha_core/n12374_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [16])
);
defparam \top/processor/sha_core/h7_16_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_15_s1  (
	.D(\top/processor/sha_core/n12375_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [15])
);
defparam \top/processor/sha_core/h7_15_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_14_s1  (
	.D(\top/processor/sha_core/n12376_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [14])
);
defparam \top/processor/sha_core/h7_14_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_13_s1  (
	.D(\top/processor/sha_core/n12377_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [13])
);
defparam \top/processor/sha_core/h7_13_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_12_s1  (
	.D(\top/processor/sha_core/n12378_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [12])
);
defparam \top/processor/sha_core/h7_12_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_11_s1  (
	.D(\top/processor/sha_core/n12379_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [11])
);
defparam \top/processor/sha_core/h7_11_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_10_s1  (
	.D(\top/processor/sha_core/n12380_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [10])
);
defparam \top/processor/sha_core/h7_10_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_9_s1  (
	.D(\top/processor/sha_core/n12381_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [9])
);
defparam \top/processor/sha_core/h7_9_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_8_s1  (
	.D(\top/processor/sha_core/n12382_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [8])
);
defparam \top/processor/sha_core/h7_8_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_7_s1  (
	.D(\top/processor/sha_core/n12383_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [7])
);
defparam \top/processor/sha_core/h7_7_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_6_s1  (
	.D(\top/processor/sha_core/n12384_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [6])
);
defparam \top/processor/sha_core/h7_6_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_5_s1  (
	.D(\top/processor/sha_core/n12385_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [5])
);
defparam \top/processor/sha_core/h7_5_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_4_s1  (
	.D(\top/processor/sha_core/n12386_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [4])
);
defparam \top/processor/sha_core/h7_4_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h7_3_s1  (
	.D(\top/processor/sha_core/n12387_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [3])
);
defparam \top/processor/sha_core/h7_3_s1 .INIT=1'b1;
DFFCE \top/processor/sha_core/h7_2_s1  (
	.D(\top/processor/sha_core/n12388_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [2])
);
defparam \top/processor/sha_core/h7_2_s1 .INIT=1'b0;
DFFCE \top/processor/sha_core/h7_1_s1  (
	.D(\top/processor/sha_core/n12389_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/h7 [1])
);
defparam \top/processor/sha_core/h7_1_s1 .INIT=1'b0;
DFFPE \top/processor/sha_core/h7_0_s1  (
	.D(\top/processor/sha_core/n12390_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h7 [0])
);
defparam \top/processor/sha_core/h7_0_s1 .INIT=1'b1;
DFFPE \top/processor/sha_core/h0_30_s1  (
	.D(\top/processor/sha_core/n12136_9 ),
	.CLK(clk),
	.CE(\top/processor/sha_core/h0_31_8 ),
	.PRESET(rst),
	.Q(\top/processor/sha_core/h0 [30])
);
defparam \top/processor/sha_core/h0_30_s1 .INIT=1'b1;
DFFC \top/processor/sha_core/state_0_s5  (
	.D(\top/processor/sha_core/n11871_15 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/state [0])
);
defparam \top/processor/sha_core/state_0_s5 .INIT=1'b0;
DFFC \top/processor/sha_core/state_1_s3  (
	.D(\top/processor/sha_core/n11870_15 ),
	.CLK(clk),
	.CLEAR(rst),
	.Q(\top/processor/sha_core/state [1])
);
defparam \top/processor/sha_core/state_1_s3 .INIT=1'b0;
ALU \top/processor/sha_core/n3924_s  (
	.I0(\top/processor/sha_core/n3552_3 ),
	.I1(\top/processor/sha_core/n3638_181 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n3924_2 ),
	.SUM(\top/processor/sha_core/n3924_1 )
);
defparam \top/processor/sha_core/n3924_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3923_s  (
	.I0(\top/processor/sha_core/n3553_3 ),
	.I1(\top/processor/sha_core/n3637_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3924_2 ),
	.COUT(\top/processor/sha_core/n3923_2 ),
	.SUM(\top/processor/sha_core/n3923_1 )
);
defparam \top/processor/sha_core/n3923_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3922_s  (
	.I0(\top/processor/sha_core/n3554_3 ),
	.I1(\top/processor/sha_core/n3636_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3923_2 ),
	.COUT(\top/processor/sha_core/n3922_2 ),
	.SUM(\top/processor/sha_core/n3922_1 )
);
defparam \top/processor/sha_core/n3922_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3921_s  (
	.I0(\top/processor/sha_core/n3555_3 ),
	.I1(\top/processor/sha_core/n3635_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3922_2 ),
	.COUT(\top/processor/sha_core/n3921_2 ),
	.SUM(\top/processor/sha_core/n3921_1 )
);
defparam \top/processor/sha_core/n3921_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3920_s  (
	.I0(\top/processor/sha_core/n3556_3 ),
	.I1(\top/processor/sha_core/n3634_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3921_2 ),
	.COUT(\top/processor/sha_core/n3920_2 ),
	.SUM(\top/processor/sha_core/n3920_1 )
);
defparam \top/processor/sha_core/n3920_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3919_s  (
	.I0(\top/processor/sha_core/n3557_3 ),
	.I1(\top/processor/sha_core/n3633_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3920_2 ),
	.COUT(\top/processor/sha_core/n3919_2 ),
	.SUM(\top/processor/sha_core/n3919_1 )
);
defparam \top/processor/sha_core/n3919_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3918_s  (
	.I0(\top/processor/sha_core/n3558_3 ),
	.I1(\top/processor/sha_core/n3632_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3919_2 ),
	.COUT(\top/processor/sha_core/n3918_2 ),
	.SUM(\top/processor/sha_core/n3918_1 )
);
defparam \top/processor/sha_core/n3918_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3917_s  (
	.I0(\top/processor/sha_core/n3559_3 ),
	.I1(\top/processor/sha_core/n3631_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3918_2 ),
	.COUT(\top/processor/sha_core/n3917_2 ),
	.SUM(\top/processor/sha_core/n3917_1 )
);
defparam \top/processor/sha_core/n3917_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3916_s  (
	.I0(\top/processor/sha_core/n3560_3 ),
	.I1(\top/processor/sha_core/n3630_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3917_2 ),
	.COUT(\top/processor/sha_core/n3916_2 ),
	.SUM(\top/processor/sha_core/n3916_1 )
);
defparam \top/processor/sha_core/n3916_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3915_s  (
	.I0(\top/processor/sha_core/n3561_3 ),
	.I1(\top/processor/sha_core/n3629_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3916_2 ),
	.COUT(\top/processor/sha_core/n3915_2 ),
	.SUM(\top/processor/sha_core/n3915_1 )
);
defparam \top/processor/sha_core/n3915_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3914_s  (
	.I0(\top/processor/sha_core/n3562_3 ),
	.I1(\top/processor/sha_core/n3628_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3915_2 ),
	.COUT(\top/processor/sha_core/n3914_2 ),
	.SUM(\top/processor/sha_core/n3914_1 )
);
defparam \top/processor/sha_core/n3914_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3913_s  (
	.I0(\top/processor/sha_core/n3563_3 ),
	.I1(\top/processor/sha_core/n3627_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3914_2 ),
	.COUT(\top/processor/sha_core/n3913_2 ),
	.SUM(\top/processor/sha_core/n3913_1 )
);
defparam \top/processor/sha_core/n3913_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3912_s  (
	.I0(\top/processor/sha_core/n3564_3 ),
	.I1(\top/processor/sha_core/n3626_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3913_2 ),
	.COUT(\top/processor/sha_core/n3912_2 ),
	.SUM(\top/processor/sha_core/n3912_1 )
);
defparam \top/processor/sha_core/n3912_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3911_s  (
	.I0(\top/processor/sha_core/n3565_3 ),
	.I1(\top/processor/sha_core/n3625_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3912_2 ),
	.COUT(\top/processor/sha_core/n3911_2 ),
	.SUM(\top/processor/sha_core/n3911_1 )
);
defparam \top/processor/sha_core/n3911_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3910_s  (
	.I0(\top/processor/sha_core/n3566_3 ),
	.I1(\top/processor/sha_core/n3624_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3911_2 ),
	.COUT(\top/processor/sha_core/n3910_2 ),
	.SUM(\top/processor/sha_core/n3910_1 )
);
defparam \top/processor/sha_core/n3910_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3909_s  (
	.I0(\top/processor/sha_core/n3567_3 ),
	.I1(\top/processor/sha_core/n3623_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3910_2 ),
	.COUT(\top/processor/sha_core/n3909_2 ),
	.SUM(\top/processor/sha_core/n3909_1 )
);
defparam \top/processor/sha_core/n3909_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3908_s  (
	.I0(\top/processor/sha_core/n3568_3 ),
	.I1(\top/processor/sha_core/n3622_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3909_2 ),
	.COUT(\top/processor/sha_core/n3908_2 ),
	.SUM(\top/processor/sha_core/n3908_1 )
);
defparam \top/processor/sha_core/n3908_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3907_s  (
	.I0(\top/processor/sha_core/n3569_3 ),
	.I1(\top/processor/sha_core/n3621_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3908_2 ),
	.COUT(\top/processor/sha_core/n3907_2 ),
	.SUM(\top/processor/sha_core/n3907_1 )
);
defparam \top/processor/sha_core/n3907_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3906_s  (
	.I0(\top/processor/sha_core/n3570_3 ),
	.I1(\top/processor/sha_core/n3620_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3907_2 ),
	.COUT(\top/processor/sha_core/n3906_2 ),
	.SUM(\top/processor/sha_core/n3906_1 )
);
defparam \top/processor/sha_core/n3906_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3905_s  (
	.I0(\top/processor/sha_core/n3571_3 ),
	.I1(\top/processor/sha_core/n3619_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3906_2 ),
	.COUT(\top/processor/sha_core/n3905_2 ),
	.SUM(\top/processor/sha_core/n3905_1 )
);
defparam \top/processor/sha_core/n3905_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3904_s  (
	.I0(\top/processor/sha_core/n3572_3 ),
	.I1(\top/processor/sha_core/n3618_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3905_2 ),
	.COUT(\top/processor/sha_core/n3904_2 ),
	.SUM(\top/processor/sha_core/n3904_1 )
);
defparam \top/processor/sha_core/n3904_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3903_s  (
	.I0(\top/processor/sha_core/n3573_3 ),
	.I1(\top/processor/sha_core/n3617_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3904_2 ),
	.COUT(\top/processor/sha_core/n3903_2 ),
	.SUM(\top/processor/sha_core/n3903_1 )
);
defparam \top/processor/sha_core/n3903_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3902_s  (
	.I0(\top/processor/sha_core/n3542_5 ),
	.I1(\top/processor/sha_core/n3616_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3903_2 ),
	.COUT(\top/processor/sha_core/n3902_2 ),
	.SUM(\top/processor/sha_core/n3902_1 )
);
defparam \top/processor/sha_core/n3902_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3901_s  (
	.I0(\top/processor/sha_core/n3543_3 ),
	.I1(\top/processor/sha_core/n3615_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3902_2 ),
	.COUT(\top/processor/sha_core/n3901_2 ),
	.SUM(\top/processor/sha_core/n3901_1 )
);
defparam \top/processor/sha_core/n3901_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3900_s  (
	.I0(\top/processor/sha_core/n3544_5 ),
	.I1(\top/processor/sha_core/n3614_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3901_2 ),
	.COUT(\top/processor/sha_core/n3900_2 ),
	.SUM(\top/processor/sha_core/n3900_1 )
);
defparam \top/processor/sha_core/n3900_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3899_s  (
	.I0(\top/processor/sha_core/n3545_3 ),
	.I1(\top/processor/sha_core/n3613_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3900_2 ),
	.COUT(\top/processor/sha_core/n3899_2 ),
	.SUM(\top/processor/sha_core/n3899_1 )
);
defparam \top/processor/sha_core/n3899_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3898_s  (
	.I0(\top/processor/sha_core/n3546_3 ),
	.I1(\top/processor/sha_core/n3612_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3899_2 ),
	.COUT(\top/processor/sha_core/n3898_2 ),
	.SUM(\top/processor/sha_core/n3898_1 )
);
defparam \top/processor/sha_core/n3898_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3897_s  (
	.I0(\top/processor/sha_core/n3547_3 ),
	.I1(\top/processor/sha_core/n3611_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3898_2 ),
	.COUT(\top/processor/sha_core/n3897_2 ),
	.SUM(\top/processor/sha_core/n3897_1 )
);
defparam \top/processor/sha_core/n3897_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3896_s  (
	.I0(\top/processor/sha_core/n3548_3 ),
	.I1(\top/processor/sha_core/n3610_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3897_2 ),
	.COUT(\top/processor/sha_core/n3896_2 ),
	.SUM(\top/processor/sha_core/n3896_1 )
);
defparam \top/processor/sha_core/n3896_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3895_s  (
	.I0(\top/processor/sha_core/n3549_3 ),
	.I1(\top/processor/sha_core/n3609_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3896_2 ),
	.COUT(\top/processor/sha_core/n3895_2 ),
	.SUM(\top/processor/sha_core/n3895_1 )
);
defparam \top/processor/sha_core/n3895_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3894_s  (
	.I0(\top/processor/sha_core/n3550_3 ),
	.I1(\top/processor/sha_core/n3608_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3895_2 ),
	.COUT(\top/processor/sha_core/n3894_2 ),
	.SUM(\top/processor/sha_core/n3894_1 )
);
defparam \top/processor/sha_core/n3894_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3893_s  (
	.I0(\top/processor/sha_core/n3551_3 ),
	.I1(\top/processor/sha_core/n3607_181 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3894_2 ),
	.COUT(\top/processor/sha_core/n3893_0_COUT ),
	.SUM(\top/processor/sha_core/n3893_1 )
);
defparam \top/processor/sha_core/n3893_s .ALU_MODE=0;
ALU \top/processor/sha_core/n3924_s0  (
	.I0(\top/processor/sha_core/n3769_3 ),
	.I1(\top/processor/sha_core/n3891_145 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n3924_4 ),
	.SUM(\top/processor/sha_core/n3924_3 )
);
defparam \top/processor/sha_core/n3924_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3923_s0  (
	.I0(\top/processor/sha_core/n3770_3 ),
	.I1(\top/processor/sha_core/n3890_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3924_4 ),
	.COUT(\top/processor/sha_core/n3923_4 ),
	.SUM(\top/processor/sha_core/n3923_3 )
);
defparam \top/processor/sha_core/n3923_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3922_s0  (
	.I0(\top/processor/sha_core/n3771_3 ),
	.I1(\top/processor/sha_core/n3889_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3923_4 ),
	.COUT(\top/processor/sha_core/n3922_4 ),
	.SUM(\top/processor/sha_core/n3922_3 )
);
defparam \top/processor/sha_core/n3922_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3921_s0  (
	.I0(\top/processor/sha_core/n3772_3 ),
	.I1(\top/processor/sha_core/n3888_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3922_4 ),
	.COUT(\top/processor/sha_core/n3921_4 ),
	.SUM(\top/processor/sha_core/n3921_3 )
);
defparam \top/processor/sha_core/n3921_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3920_s0  (
	.I0(\top/processor/sha_core/n3773_3 ),
	.I1(\top/processor/sha_core/n3887_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3921_4 ),
	.COUT(\top/processor/sha_core/n3920_4 ),
	.SUM(\top/processor/sha_core/n3920_3 )
);
defparam \top/processor/sha_core/n3920_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3919_s0  (
	.I0(\top/processor/sha_core/n3774_3 ),
	.I1(\top/processor/sha_core/n3886_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3920_4 ),
	.COUT(\top/processor/sha_core/n3919_4 ),
	.SUM(\top/processor/sha_core/n3919_3 )
);
defparam \top/processor/sha_core/n3919_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3918_s0  (
	.I0(\top/processor/sha_core/n3775_3 ),
	.I1(\top/processor/sha_core/n3885_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3919_4 ),
	.COUT(\top/processor/sha_core/n3918_4 ),
	.SUM(\top/processor/sha_core/n3918_3 )
);
defparam \top/processor/sha_core/n3918_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3917_s0  (
	.I0(\top/processor/sha_core/n3776_3 ),
	.I1(\top/processor/sha_core/n3884_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3918_4 ),
	.COUT(\top/processor/sha_core/n3917_4 ),
	.SUM(\top/processor/sha_core/n3917_3 )
);
defparam \top/processor/sha_core/n3917_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3916_s0  (
	.I0(\top/processor/sha_core/n3777_3 ),
	.I1(\top/processor/sha_core/n3883_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3917_4 ),
	.COUT(\top/processor/sha_core/n3916_4 ),
	.SUM(\top/processor/sha_core/n3916_3 )
);
defparam \top/processor/sha_core/n3916_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3915_s0  (
	.I0(\top/processor/sha_core/n3778_3 ),
	.I1(\top/processor/sha_core/n3882_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3916_4 ),
	.COUT(\top/processor/sha_core/n3915_4 ),
	.SUM(\top/processor/sha_core/n3915_3 )
);
defparam \top/processor/sha_core/n3915_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3914_s0  (
	.I0(\top/processor/sha_core/n3779_3 ),
	.I1(\top/processor/sha_core/n3881_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3915_4 ),
	.COUT(\top/processor/sha_core/n3914_4 ),
	.SUM(\top/processor/sha_core/n3914_3 )
);
defparam \top/processor/sha_core/n3914_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3913_s0  (
	.I0(\top/processor/sha_core/n3780_3 ),
	.I1(\top/processor/sha_core/n3880_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3914_4 ),
	.COUT(\top/processor/sha_core/n3913_4 ),
	.SUM(\top/processor/sha_core/n3913_3 )
);
defparam \top/processor/sha_core/n3913_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3912_s0  (
	.I0(\top/processor/sha_core/n3781_3 ),
	.I1(\top/processor/sha_core/n3879_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3913_4 ),
	.COUT(\top/processor/sha_core/n3912_4 ),
	.SUM(\top/processor/sha_core/n3912_3 )
);
defparam \top/processor/sha_core/n3912_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3911_s0  (
	.I0(\top/processor/sha_core/n3782_3 ),
	.I1(\top/processor/sha_core/n3878_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3912_4 ),
	.COUT(\top/processor/sha_core/n3911_4 ),
	.SUM(\top/processor/sha_core/n3911_3 )
);
defparam \top/processor/sha_core/n3911_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3910_s0  (
	.I0(\top/processor/sha_core/n3783_3 ),
	.I1(\top/processor/sha_core/n3877_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3911_4 ),
	.COUT(\top/processor/sha_core/n3910_4 ),
	.SUM(\top/processor/sha_core/n3910_3 )
);
defparam \top/processor/sha_core/n3910_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3909_s0  (
	.I0(\top/processor/sha_core/n3784_3 ),
	.I1(\top/processor/sha_core/n3876_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3910_4 ),
	.COUT(\top/processor/sha_core/n3909_4 ),
	.SUM(\top/processor/sha_core/n3909_3 )
);
defparam \top/processor/sha_core/n3909_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3908_s0  (
	.I0(\top/processor/sha_core/n3785_3 ),
	.I1(\top/processor/sha_core/n3875_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3909_4 ),
	.COUT(\top/processor/sha_core/n3908_4 ),
	.SUM(\top/processor/sha_core/n3908_3 )
);
defparam \top/processor/sha_core/n3908_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3907_s0  (
	.I0(\top/processor/sha_core/n3786_3 ),
	.I1(\top/processor/sha_core/n3874_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3908_4 ),
	.COUT(\top/processor/sha_core/n3907_4 ),
	.SUM(\top/processor/sha_core/n3907_3 )
);
defparam \top/processor/sha_core/n3907_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3906_s0  (
	.I0(\top/processor/sha_core/n3787_3 ),
	.I1(\top/processor/sha_core/n3873_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3907_4 ),
	.COUT(\top/processor/sha_core/n3906_4 ),
	.SUM(\top/processor/sha_core/n3906_3 )
);
defparam \top/processor/sha_core/n3906_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3905_s0  (
	.I0(\top/processor/sha_core/n3788_3 ),
	.I1(\top/processor/sha_core/n3872_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3906_4 ),
	.COUT(\top/processor/sha_core/n3905_4 ),
	.SUM(\top/processor/sha_core/n3905_3 )
);
defparam \top/processor/sha_core/n3905_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3904_s0  (
	.I0(\top/processor/sha_core/n3789_3 ),
	.I1(\top/processor/sha_core/n3871_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3905_4 ),
	.COUT(\top/processor/sha_core/n3904_4 ),
	.SUM(\top/processor/sha_core/n3904_3 )
);
defparam \top/processor/sha_core/n3904_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3903_s0  (
	.I0(\top/processor/sha_core/n3790_3 ),
	.I1(\top/processor/sha_core/n3870_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3904_4 ),
	.COUT(\top/processor/sha_core/n3903_4 ),
	.SUM(\top/processor/sha_core/n3903_3 )
);
defparam \top/processor/sha_core/n3903_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3902_s0  (
	.I0(\top/processor/sha_core/n3791_3 ),
	.I1(\top/processor/sha_core/n3869_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3903_4 ),
	.COUT(\top/processor/sha_core/n3902_4 ),
	.SUM(\top/processor/sha_core/n3902_3 )
);
defparam \top/processor/sha_core/n3902_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3901_s0  (
	.I0(\top/processor/sha_core/n3792_3 ),
	.I1(\top/processor/sha_core/n3868_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3902_4 ),
	.COUT(\top/processor/sha_core/n3901_4 ),
	.SUM(\top/processor/sha_core/n3901_3 )
);
defparam \top/processor/sha_core/n3901_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3900_s0  (
	.I0(\top/processor/sha_core/n3793_3 ),
	.I1(\top/processor/sha_core/n3867_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3901_4 ),
	.COUT(\top/processor/sha_core/n3900_4 ),
	.SUM(\top/processor/sha_core/n3900_3 )
);
defparam \top/processor/sha_core/n3900_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3899_s0  (
	.I0(\top/processor/sha_core/n3794_3 ),
	.I1(\top/processor/sha_core/n3866_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3900_4 ),
	.COUT(\top/processor/sha_core/n3899_4 ),
	.SUM(\top/processor/sha_core/n3899_3 )
);
defparam \top/processor/sha_core/n3899_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3898_s0  (
	.I0(\top/processor/sha_core/n3795_3 ),
	.I1(\top/processor/sha_core/n3865_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3899_4 ),
	.COUT(\top/processor/sha_core/n3898_4 ),
	.SUM(\top/processor/sha_core/n3898_3 )
);
defparam \top/processor/sha_core/n3898_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3897_s0  (
	.I0(\top/processor/sha_core/n3796_3 ),
	.I1(\top/processor/sha_core/n3864_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3898_4 ),
	.COUT(\top/processor/sha_core/n3897_4 ),
	.SUM(\top/processor/sha_core/n3897_3 )
);
defparam \top/processor/sha_core/n3897_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3896_s0  (
	.I0(\top/processor/sha_core/n3797_3 ),
	.I1(\top/processor/sha_core/n3863_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3897_4 ),
	.COUT(\top/processor/sha_core/n3896_4 ),
	.SUM(\top/processor/sha_core/n3896_3 )
);
defparam \top/processor/sha_core/n3896_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3895_s0  (
	.I0(\top/processor/sha_core/n3766_16 ),
	.I1(\top/processor/sha_core/n3862_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3896_4 ),
	.COUT(\top/processor/sha_core/n3895_4 ),
	.SUM(\top/processor/sha_core/n3895_3 )
);
defparam \top/processor/sha_core/n3895_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3894_s0  (
	.I0(\top/processor/sha_core/n3767_15 ),
	.I1(\top/processor/sha_core/n3861_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3895_4 ),
	.COUT(\top/processor/sha_core/n3894_4 ),
	.SUM(\top/processor/sha_core/n3894_3 )
);
defparam \top/processor/sha_core/n3894_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3893_s0  (
	.I0(\top/processor/sha_core/n3768_15 ),
	.I1(\top/processor/sha_core/n3860_145 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3894_4 ),
	.COUT(\top/processor/sha_core/n3893_1_COUT ),
	.SUM(\top/processor/sha_core/n3893_3 )
);
defparam \top/processor/sha_core/n3893_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n3924_s1  (
	.I0(\top/processor/sha_core/n3924_1 ),
	.I1(\top/processor/sha_core/n3924_3 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n3924_6 ),
	.SUM(\top/processor/sha_core/n3924_5 )
);
defparam \top/processor/sha_core/n3924_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3923_s1  (
	.I0(\top/processor/sha_core/n3923_1 ),
	.I1(\top/processor/sha_core/n3923_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3924_6 ),
	.COUT(\top/processor/sha_core/n3923_6 ),
	.SUM(\top/processor/sha_core/n3923_5 )
);
defparam \top/processor/sha_core/n3923_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3922_s1  (
	.I0(\top/processor/sha_core/n3922_1 ),
	.I1(\top/processor/sha_core/n3922_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3923_6 ),
	.COUT(\top/processor/sha_core/n3922_6 ),
	.SUM(\top/processor/sha_core/n3922_5 )
);
defparam \top/processor/sha_core/n3922_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3921_s1  (
	.I0(\top/processor/sha_core/n3921_1 ),
	.I1(\top/processor/sha_core/n3921_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3922_6 ),
	.COUT(\top/processor/sha_core/n3921_6 ),
	.SUM(\top/processor/sha_core/n3921_5 )
);
defparam \top/processor/sha_core/n3921_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3920_s1  (
	.I0(\top/processor/sha_core/n3920_1 ),
	.I1(\top/processor/sha_core/n3920_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3921_6 ),
	.COUT(\top/processor/sha_core/n3920_6 ),
	.SUM(\top/processor/sha_core/n3920_5 )
);
defparam \top/processor/sha_core/n3920_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3919_s1  (
	.I0(\top/processor/sha_core/n3919_1 ),
	.I1(\top/processor/sha_core/n3919_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3920_6 ),
	.COUT(\top/processor/sha_core/n3919_6 ),
	.SUM(\top/processor/sha_core/n3919_5 )
);
defparam \top/processor/sha_core/n3919_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3918_s1  (
	.I0(\top/processor/sha_core/n3918_1 ),
	.I1(\top/processor/sha_core/n3918_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3919_6 ),
	.COUT(\top/processor/sha_core/n3918_6 ),
	.SUM(\top/processor/sha_core/n3918_5 )
);
defparam \top/processor/sha_core/n3918_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3917_s1  (
	.I0(\top/processor/sha_core/n3917_1 ),
	.I1(\top/processor/sha_core/n3917_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3918_6 ),
	.COUT(\top/processor/sha_core/n3917_6 ),
	.SUM(\top/processor/sha_core/n3917_5 )
);
defparam \top/processor/sha_core/n3917_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3916_s1  (
	.I0(\top/processor/sha_core/n3916_1 ),
	.I1(\top/processor/sha_core/n3916_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3917_6 ),
	.COUT(\top/processor/sha_core/n3916_6 ),
	.SUM(\top/processor/sha_core/n3916_5 )
);
defparam \top/processor/sha_core/n3916_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3915_s1  (
	.I0(\top/processor/sha_core/n3915_1 ),
	.I1(\top/processor/sha_core/n3915_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3916_6 ),
	.COUT(\top/processor/sha_core/n3915_6 ),
	.SUM(\top/processor/sha_core/n3915_5 )
);
defparam \top/processor/sha_core/n3915_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3914_s1  (
	.I0(\top/processor/sha_core/n3914_1 ),
	.I1(\top/processor/sha_core/n3914_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3915_6 ),
	.COUT(\top/processor/sha_core/n3914_6 ),
	.SUM(\top/processor/sha_core/n3914_5 )
);
defparam \top/processor/sha_core/n3914_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3913_s1  (
	.I0(\top/processor/sha_core/n3913_1 ),
	.I1(\top/processor/sha_core/n3913_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3914_6 ),
	.COUT(\top/processor/sha_core/n3913_6 ),
	.SUM(\top/processor/sha_core/n3913_5 )
);
defparam \top/processor/sha_core/n3913_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3912_s1  (
	.I0(\top/processor/sha_core/n3912_1 ),
	.I1(\top/processor/sha_core/n3912_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3913_6 ),
	.COUT(\top/processor/sha_core/n3912_6 ),
	.SUM(\top/processor/sha_core/n3912_5 )
);
defparam \top/processor/sha_core/n3912_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3911_s1  (
	.I0(\top/processor/sha_core/n3911_1 ),
	.I1(\top/processor/sha_core/n3911_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3912_6 ),
	.COUT(\top/processor/sha_core/n3911_6 ),
	.SUM(\top/processor/sha_core/n3911_5 )
);
defparam \top/processor/sha_core/n3911_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3910_s1  (
	.I0(\top/processor/sha_core/n3910_1 ),
	.I1(\top/processor/sha_core/n3910_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3911_6 ),
	.COUT(\top/processor/sha_core/n3910_6 ),
	.SUM(\top/processor/sha_core/n3910_5 )
);
defparam \top/processor/sha_core/n3910_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3909_s1  (
	.I0(\top/processor/sha_core/n3909_1 ),
	.I1(\top/processor/sha_core/n3909_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3910_6 ),
	.COUT(\top/processor/sha_core/n3909_6 ),
	.SUM(\top/processor/sha_core/n3909_5 )
);
defparam \top/processor/sha_core/n3909_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3908_s1  (
	.I0(\top/processor/sha_core/n3908_1 ),
	.I1(\top/processor/sha_core/n3908_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3909_6 ),
	.COUT(\top/processor/sha_core/n3908_6 ),
	.SUM(\top/processor/sha_core/n3908_5 )
);
defparam \top/processor/sha_core/n3908_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3907_s1  (
	.I0(\top/processor/sha_core/n3907_1 ),
	.I1(\top/processor/sha_core/n3907_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3908_6 ),
	.COUT(\top/processor/sha_core/n3907_6 ),
	.SUM(\top/processor/sha_core/n3907_5 )
);
defparam \top/processor/sha_core/n3907_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3906_s1  (
	.I0(\top/processor/sha_core/n3906_1 ),
	.I1(\top/processor/sha_core/n3906_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3907_6 ),
	.COUT(\top/processor/sha_core/n3906_6 ),
	.SUM(\top/processor/sha_core/n3906_5 )
);
defparam \top/processor/sha_core/n3906_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3905_s1  (
	.I0(\top/processor/sha_core/n3905_1 ),
	.I1(\top/processor/sha_core/n3905_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3906_6 ),
	.COUT(\top/processor/sha_core/n3905_6 ),
	.SUM(\top/processor/sha_core/n3905_5 )
);
defparam \top/processor/sha_core/n3905_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3904_s1  (
	.I0(\top/processor/sha_core/n3904_1 ),
	.I1(\top/processor/sha_core/n3904_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3905_6 ),
	.COUT(\top/processor/sha_core/n3904_6 ),
	.SUM(\top/processor/sha_core/n3904_5 )
);
defparam \top/processor/sha_core/n3904_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3903_s1  (
	.I0(\top/processor/sha_core/n3903_1 ),
	.I1(\top/processor/sha_core/n3903_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3904_6 ),
	.COUT(\top/processor/sha_core/n3903_6 ),
	.SUM(\top/processor/sha_core/n3903_5 )
);
defparam \top/processor/sha_core/n3903_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3902_s1  (
	.I0(\top/processor/sha_core/n3902_1 ),
	.I1(\top/processor/sha_core/n3902_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3903_6 ),
	.COUT(\top/processor/sha_core/n3902_6 ),
	.SUM(\top/processor/sha_core/n3902_5 )
);
defparam \top/processor/sha_core/n3902_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3901_s1  (
	.I0(\top/processor/sha_core/n3901_1 ),
	.I1(\top/processor/sha_core/n3901_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3902_6 ),
	.COUT(\top/processor/sha_core/n3901_6 ),
	.SUM(\top/processor/sha_core/n3901_5 )
);
defparam \top/processor/sha_core/n3901_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3900_s1  (
	.I0(\top/processor/sha_core/n3900_1 ),
	.I1(\top/processor/sha_core/n3900_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3901_6 ),
	.COUT(\top/processor/sha_core/n3900_6 ),
	.SUM(\top/processor/sha_core/n3900_5 )
);
defparam \top/processor/sha_core/n3900_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3899_s1  (
	.I0(\top/processor/sha_core/n3899_1 ),
	.I1(\top/processor/sha_core/n3899_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3900_6 ),
	.COUT(\top/processor/sha_core/n3899_6 ),
	.SUM(\top/processor/sha_core/n3899_5 )
);
defparam \top/processor/sha_core/n3899_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3898_s1  (
	.I0(\top/processor/sha_core/n3898_1 ),
	.I1(\top/processor/sha_core/n3898_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3899_6 ),
	.COUT(\top/processor/sha_core/n3898_6 ),
	.SUM(\top/processor/sha_core/n3898_5 )
);
defparam \top/processor/sha_core/n3898_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3897_s1  (
	.I0(\top/processor/sha_core/n3897_1 ),
	.I1(\top/processor/sha_core/n3897_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3898_6 ),
	.COUT(\top/processor/sha_core/n3897_6 ),
	.SUM(\top/processor/sha_core/n3897_5 )
);
defparam \top/processor/sha_core/n3897_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3896_s1  (
	.I0(\top/processor/sha_core/n3896_1 ),
	.I1(\top/processor/sha_core/n3896_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3897_6 ),
	.COUT(\top/processor/sha_core/n3896_6 ),
	.SUM(\top/processor/sha_core/n3896_5 )
);
defparam \top/processor/sha_core/n3896_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3895_s1  (
	.I0(\top/processor/sha_core/n3895_1 ),
	.I1(\top/processor/sha_core/n3895_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3896_6 ),
	.COUT(\top/processor/sha_core/n3895_6 ),
	.SUM(\top/processor/sha_core/n3895_5 )
);
defparam \top/processor/sha_core/n3895_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3894_s1  (
	.I0(\top/processor/sha_core/n3894_1 ),
	.I1(\top/processor/sha_core/n3894_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3895_6 ),
	.COUT(\top/processor/sha_core/n3894_6 ),
	.SUM(\top/processor/sha_core/n3894_5 )
);
defparam \top/processor/sha_core/n3894_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n3893_s1  (
	.I0(\top/processor/sha_core/n3893_1 ),
	.I1(\top/processor/sha_core/n3893_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n3894_6 ),
	.COUT(\top/processor/sha_core/n3893_2_COUT ),
	.SUM(\top/processor/sha_core/n3893_5 )
);
defparam \top/processor/sha_core/n3893_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10857_s  (
	.I0(\top/processor/sha_core/h0 [0]),
	.I1(\top/processor/sha_core/a [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10857_2 ),
	.SUM(\top/processor/sha_core/n10857_1 )
);
defparam \top/processor/sha_core/n10857_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10856_s  (
	.I0(\top/processor/sha_core/h0 [1]),
	.I1(\top/processor/sha_core/a [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10857_2 ),
	.COUT(\top/processor/sha_core/n10856_2 ),
	.SUM(\top/processor/sha_core/n10856_1 )
);
defparam \top/processor/sha_core/n10856_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10855_s  (
	.I0(\top/processor/sha_core/h0 [2]),
	.I1(\top/processor/sha_core/a [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10856_2 ),
	.COUT(\top/processor/sha_core/n10855_2 ),
	.SUM(\top/processor/sha_core/n10855_1 )
);
defparam \top/processor/sha_core/n10855_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10854_s  (
	.I0(\top/processor/sha_core/h0 [3]),
	.I1(\top/processor/sha_core/a [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10855_2 ),
	.COUT(\top/processor/sha_core/n10854_2 ),
	.SUM(\top/processor/sha_core/n10854_1 )
);
defparam \top/processor/sha_core/n10854_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10853_s  (
	.I0(\top/processor/sha_core/h0 [4]),
	.I1(\top/processor/sha_core/a [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10854_2 ),
	.COUT(\top/processor/sha_core/n10853_2 ),
	.SUM(\top/processor/sha_core/n10853_1 )
);
defparam \top/processor/sha_core/n10853_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10852_s  (
	.I0(\top/processor/sha_core/h0 [5]),
	.I1(\top/processor/sha_core/a [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10853_2 ),
	.COUT(\top/processor/sha_core/n10852_2 ),
	.SUM(\top/processor/sha_core/n10852_1 )
);
defparam \top/processor/sha_core/n10852_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10851_s  (
	.I0(\top/processor/sha_core/h0 [6]),
	.I1(\top/processor/sha_core/a [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10852_2 ),
	.COUT(\top/processor/sha_core/n10851_2 ),
	.SUM(\top/processor/sha_core/n10851_1 )
);
defparam \top/processor/sha_core/n10851_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10850_s  (
	.I0(\top/processor/sha_core/h0 [7]),
	.I1(\top/processor/sha_core/a [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10851_2 ),
	.COUT(\top/processor/sha_core/n10850_2 ),
	.SUM(\top/processor/sha_core/n10850_1 )
);
defparam \top/processor/sha_core/n10850_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10849_s  (
	.I0(\top/processor/sha_core/h0 [8]),
	.I1(\top/processor/sha_core/a [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10850_2 ),
	.COUT(\top/processor/sha_core/n10849_2 ),
	.SUM(\top/processor/sha_core/n10849_1 )
);
defparam \top/processor/sha_core/n10849_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10848_s  (
	.I0(\top/processor/sha_core/h0 [9]),
	.I1(\top/processor/sha_core/a [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10849_2 ),
	.COUT(\top/processor/sha_core/n10848_2 ),
	.SUM(\top/processor/sha_core/n10848_1 )
);
defparam \top/processor/sha_core/n10848_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10847_s  (
	.I0(\top/processor/sha_core/h0 [10]),
	.I1(\top/processor/sha_core/a [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10848_2 ),
	.COUT(\top/processor/sha_core/n10847_2 ),
	.SUM(\top/processor/sha_core/n10847_1 )
);
defparam \top/processor/sha_core/n10847_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10846_s  (
	.I0(\top/processor/sha_core/h0 [11]),
	.I1(\top/processor/sha_core/a [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10847_2 ),
	.COUT(\top/processor/sha_core/n10846_2 ),
	.SUM(\top/processor/sha_core/n10846_1 )
);
defparam \top/processor/sha_core/n10846_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10845_s  (
	.I0(\top/processor/sha_core/h0 [12]),
	.I1(\top/processor/sha_core/a [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10846_2 ),
	.COUT(\top/processor/sha_core/n10845_2 ),
	.SUM(\top/processor/sha_core/n10845_1 )
);
defparam \top/processor/sha_core/n10845_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10844_s  (
	.I0(\top/processor/sha_core/h0 [13]),
	.I1(\top/processor/sha_core/a [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10845_2 ),
	.COUT(\top/processor/sha_core/n10844_2 ),
	.SUM(\top/processor/sha_core/n10844_1 )
);
defparam \top/processor/sha_core/n10844_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10843_s  (
	.I0(\top/processor/sha_core/h0 [14]),
	.I1(\top/processor/sha_core/a [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10844_2 ),
	.COUT(\top/processor/sha_core/n10843_2 ),
	.SUM(\top/processor/sha_core/n10843_1 )
);
defparam \top/processor/sha_core/n10843_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10842_s  (
	.I0(\top/processor/sha_core/h0 [15]),
	.I1(\top/processor/sha_core/a [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10843_2 ),
	.COUT(\top/processor/sha_core/n10842_2 ),
	.SUM(\top/processor/sha_core/n10842_1 )
);
defparam \top/processor/sha_core/n10842_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10841_s  (
	.I0(\top/processor/sha_core/h0 [16]),
	.I1(\top/processor/sha_core/a [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10842_2 ),
	.COUT(\top/processor/sha_core/n10841_2 ),
	.SUM(\top/processor/sha_core/n10841_1 )
);
defparam \top/processor/sha_core/n10841_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10840_s  (
	.I0(\top/processor/sha_core/h0 [17]),
	.I1(\top/processor/sha_core/a [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10841_2 ),
	.COUT(\top/processor/sha_core/n10840_2 ),
	.SUM(\top/processor/sha_core/n10840_1 )
);
defparam \top/processor/sha_core/n10840_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10839_s  (
	.I0(\top/processor/sha_core/h0 [18]),
	.I1(\top/processor/sha_core/a [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10840_2 ),
	.COUT(\top/processor/sha_core/n10839_2 ),
	.SUM(\top/processor/sha_core/n10839_1 )
);
defparam \top/processor/sha_core/n10839_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10838_s  (
	.I0(\top/processor/sha_core/h0 [19]),
	.I1(\top/processor/sha_core/a [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10839_2 ),
	.COUT(\top/processor/sha_core/n10838_2 ),
	.SUM(\top/processor/sha_core/n10838_1 )
);
defparam \top/processor/sha_core/n10838_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10837_s  (
	.I0(\top/processor/sha_core/h0 [20]),
	.I1(\top/processor/sha_core/a [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10838_2 ),
	.COUT(\top/processor/sha_core/n10837_2 ),
	.SUM(\top/processor/sha_core/n10837_1 )
);
defparam \top/processor/sha_core/n10837_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10836_s  (
	.I0(\top/processor/sha_core/h0 [21]),
	.I1(\top/processor/sha_core/a [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10837_2 ),
	.COUT(\top/processor/sha_core/n10836_2 ),
	.SUM(\top/processor/sha_core/n10836_1 )
);
defparam \top/processor/sha_core/n10836_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10835_s  (
	.I0(\top/processor/sha_core/h0 [22]),
	.I1(\top/processor/sha_core/a [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10836_2 ),
	.COUT(\top/processor/sha_core/n10835_2 ),
	.SUM(\top/processor/sha_core/n10835_1 )
);
defparam \top/processor/sha_core/n10835_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10834_s  (
	.I0(\top/processor/sha_core/h0 [23]),
	.I1(\top/processor/sha_core/a [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10835_2 ),
	.COUT(\top/processor/sha_core/n10834_2 ),
	.SUM(\top/processor/sha_core/n10834_1 )
);
defparam \top/processor/sha_core/n10834_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10833_s  (
	.I0(\top/processor/sha_core/h0 [24]),
	.I1(\top/processor/sha_core/a [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10834_2 ),
	.COUT(\top/processor/sha_core/n10833_2 ),
	.SUM(\top/processor/sha_core/n10833_1 )
);
defparam \top/processor/sha_core/n10833_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10832_s  (
	.I0(\top/processor/sha_core/h0 [25]),
	.I1(\top/processor/sha_core/a [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10833_2 ),
	.COUT(\top/processor/sha_core/n10832_2 ),
	.SUM(\top/processor/sha_core/n10832_1 )
);
defparam \top/processor/sha_core/n10832_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10831_s  (
	.I0(\top/processor/sha_core/h0 [26]),
	.I1(\top/processor/sha_core/a [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10832_2 ),
	.COUT(\top/processor/sha_core/n10831_2 ),
	.SUM(\top/processor/sha_core/n10831_1 )
);
defparam \top/processor/sha_core/n10831_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10830_s  (
	.I0(\top/processor/sha_core/h0 [27]),
	.I1(\top/processor/sha_core/a [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10831_2 ),
	.COUT(\top/processor/sha_core/n10830_2 ),
	.SUM(\top/processor/sha_core/n10830_1 )
);
defparam \top/processor/sha_core/n10830_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10829_s  (
	.I0(\top/processor/sha_core/h0 [28]),
	.I1(\top/processor/sha_core/a [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10830_2 ),
	.COUT(\top/processor/sha_core/n10829_2 ),
	.SUM(\top/processor/sha_core/n10829_1 )
);
defparam \top/processor/sha_core/n10829_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10828_s  (
	.I0(\top/processor/sha_core/h0 [29]),
	.I1(\top/processor/sha_core/a [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10829_2 ),
	.COUT(\top/processor/sha_core/n10828_2 ),
	.SUM(\top/processor/sha_core/n10828_1 )
);
defparam \top/processor/sha_core/n10828_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10827_s  (
	.I0(\top/processor/sha_core/h0 [30]),
	.I1(\top/processor/sha_core/a [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10828_2 ),
	.COUT(\top/processor/sha_core/n10827_2 ),
	.SUM(\top/processor/sha_core/n10827_1 )
);
defparam \top/processor/sha_core/n10827_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10826_s  (
	.I0(\top/processor/sha_core/h0 [31]),
	.I1(\top/processor/sha_core/a [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10827_2 ),
	.COUT(\top/processor/sha_core/n10826_0_COUT ),
	.SUM(\top/processor/sha_core/n10826_1 )
);
defparam \top/processor/sha_core/n10826_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10890_s  (
	.I0(\top/processor/sha_core/h1 [0]),
	.I1(\top/processor/sha_core/b [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10890_2 ),
	.SUM(\top/processor/sha_core/n10890_1 )
);
defparam \top/processor/sha_core/n10890_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10889_s  (
	.I0(\top/processor/sha_core/h1 [1]),
	.I1(\top/processor/sha_core/b [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10890_2 ),
	.COUT(\top/processor/sha_core/n10889_2 ),
	.SUM(\top/processor/sha_core/n10889_1 )
);
defparam \top/processor/sha_core/n10889_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10888_s  (
	.I0(\top/processor/sha_core/h1 [2]),
	.I1(\top/processor/sha_core/b [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10889_2 ),
	.COUT(\top/processor/sha_core/n10888_2 ),
	.SUM(\top/processor/sha_core/n10888_1 )
);
defparam \top/processor/sha_core/n10888_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10887_s  (
	.I0(\top/processor/sha_core/h1 [3]),
	.I1(\top/processor/sha_core/b [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10888_2 ),
	.COUT(\top/processor/sha_core/n10887_2 ),
	.SUM(\top/processor/sha_core/n10887_1 )
);
defparam \top/processor/sha_core/n10887_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10886_s  (
	.I0(\top/processor/sha_core/h1 [4]),
	.I1(\top/processor/sha_core/b [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10887_2 ),
	.COUT(\top/processor/sha_core/n10886_2 ),
	.SUM(\top/processor/sha_core/n10886_1 )
);
defparam \top/processor/sha_core/n10886_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10885_s  (
	.I0(\top/processor/sha_core/h1 [5]),
	.I1(\top/processor/sha_core/b [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10886_2 ),
	.COUT(\top/processor/sha_core/n10885_2 ),
	.SUM(\top/processor/sha_core/n10885_1 )
);
defparam \top/processor/sha_core/n10885_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10884_s  (
	.I0(\top/processor/sha_core/h1 [6]),
	.I1(\top/processor/sha_core/b [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10885_2 ),
	.COUT(\top/processor/sha_core/n10884_2 ),
	.SUM(\top/processor/sha_core/n10884_1 )
);
defparam \top/processor/sha_core/n10884_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10883_s  (
	.I0(\top/processor/sha_core/h1 [7]),
	.I1(\top/processor/sha_core/b [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10884_2 ),
	.COUT(\top/processor/sha_core/n10883_2 ),
	.SUM(\top/processor/sha_core/n10883_1 )
);
defparam \top/processor/sha_core/n10883_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10882_s  (
	.I0(\top/processor/sha_core/h1 [8]),
	.I1(\top/processor/sha_core/b [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10883_2 ),
	.COUT(\top/processor/sha_core/n10882_2 ),
	.SUM(\top/processor/sha_core/n10882_1 )
);
defparam \top/processor/sha_core/n10882_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10881_s  (
	.I0(\top/processor/sha_core/h1 [9]),
	.I1(\top/processor/sha_core/b [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10882_2 ),
	.COUT(\top/processor/sha_core/n10881_2 ),
	.SUM(\top/processor/sha_core/n10881_1 )
);
defparam \top/processor/sha_core/n10881_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10880_s  (
	.I0(\top/processor/sha_core/h1 [10]),
	.I1(\top/processor/sha_core/b [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10881_2 ),
	.COUT(\top/processor/sha_core/n10880_2 ),
	.SUM(\top/processor/sha_core/n10880_1 )
);
defparam \top/processor/sha_core/n10880_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10879_s  (
	.I0(\top/processor/sha_core/h1 [11]),
	.I1(\top/processor/sha_core/b [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10880_2 ),
	.COUT(\top/processor/sha_core/n10879_2 ),
	.SUM(\top/processor/sha_core/n10879_1 )
);
defparam \top/processor/sha_core/n10879_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10878_s  (
	.I0(\top/processor/sha_core/h1 [12]),
	.I1(\top/processor/sha_core/b [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10879_2 ),
	.COUT(\top/processor/sha_core/n10878_2 ),
	.SUM(\top/processor/sha_core/n10878_1 )
);
defparam \top/processor/sha_core/n10878_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10877_s  (
	.I0(\top/processor/sha_core/h1 [13]),
	.I1(\top/processor/sha_core/b [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10878_2 ),
	.COUT(\top/processor/sha_core/n10877_2 ),
	.SUM(\top/processor/sha_core/n10877_1 )
);
defparam \top/processor/sha_core/n10877_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10876_s  (
	.I0(\top/processor/sha_core/h1 [14]),
	.I1(\top/processor/sha_core/b [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10877_2 ),
	.COUT(\top/processor/sha_core/n10876_2 ),
	.SUM(\top/processor/sha_core/n10876_1 )
);
defparam \top/processor/sha_core/n10876_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10875_s  (
	.I0(\top/processor/sha_core/h1 [15]),
	.I1(\top/processor/sha_core/b [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10876_2 ),
	.COUT(\top/processor/sha_core/n10875_2 ),
	.SUM(\top/processor/sha_core/n10875_1 )
);
defparam \top/processor/sha_core/n10875_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10874_s  (
	.I0(\top/processor/sha_core/h1 [16]),
	.I1(\top/processor/sha_core/b [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10875_2 ),
	.COUT(\top/processor/sha_core/n10874_2 ),
	.SUM(\top/processor/sha_core/n10874_1 )
);
defparam \top/processor/sha_core/n10874_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10873_s  (
	.I0(\top/processor/sha_core/h1 [17]),
	.I1(\top/processor/sha_core/b [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10874_2 ),
	.COUT(\top/processor/sha_core/n10873_2 ),
	.SUM(\top/processor/sha_core/n10873_1 )
);
defparam \top/processor/sha_core/n10873_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10872_s  (
	.I0(\top/processor/sha_core/h1 [18]),
	.I1(\top/processor/sha_core/b [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10873_2 ),
	.COUT(\top/processor/sha_core/n10872_2 ),
	.SUM(\top/processor/sha_core/n10872_1 )
);
defparam \top/processor/sha_core/n10872_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10871_s  (
	.I0(\top/processor/sha_core/h1 [19]),
	.I1(\top/processor/sha_core/b [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10872_2 ),
	.COUT(\top/processor/sha_core/n10871_2 ),
	.SUM(\top/processor/sha_core/n10871_1 )
);
defparam \top/processor/sha_core/n10871_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10870_s  (
	.I0(\top/processor/sha_core/h1 [20]),
	.I1(\top/processor/sha_core/b [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10871_2 ),
	.COUT(\top/processor/sha_core/n10870_2 ),
	.SUM(\top/processor/sha_core/n10870_1 )
);
defparam \top/processor/sha_core/n10870_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10869_s  (
	.I0(\top/processor/sha_core/h1 [21]),
	.I1(\top/processor/sha_core/b [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10870_2 ),
	.COUT(\top/processor/sha_core/n10869_2 ),
	.SUM(\top/processor/sha_core/n10869_1 )
);
defparam \top/processor/sha_core/n10869_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10868_s  (
	.I0(\top/processor/sha_core/h1 [22]),
	.I1(\top/processor/sha_core/b [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10869_2 ),
	.COUT(\top/processor/sha_core/n10868_2 ),
	.SUM(\top/processor/sha_core/n10868_1 )
);
defparam \top/processor/sha_core/n10868_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10867_s  (
	.I0(\top/processor/sha_core/h1 [23]),
	.I1(\top/processor/sha_core/b [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10868_2 ),
	.COUT(\top/processor/sha_core/n10867_2 ),
	.SUM(\top/processor/sha_core/n10867_1 )
);
defparam \top/processor/sha_core/n10867_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10866_s  (
	.I0(\top/processor/sha_core/h1 [24]),
	.I1(\top/processor/sha_core/b [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10867_2 ),
	.COUT(\top/processor/sha_core/n10866_2 ),
	.SUM(\top/processor/sha_core/n10866_1 )
);
defparam \top/processor/sha_core/n10866_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10865_s  (
	.I0(\top/processor/sha_core/h1 [25]),
	.I1(\top/processor/sha_core/b [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10866_2 ),
	.COUT(\top/processor/sha_core/n10865_2 ),
	.SUM(\top/processor/sha_core/n10865_1 )
);
defparam \top/processor/sha_core/n10865_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10864_s  (
	.I0(\top/processor/sha_core/h1 [26]),
	.I1(\top/processor/sha_core/b [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10865_2 ),
	.COUT(\top/processor/sha_core/n10864_2 ),
	.SUM(\top/processor/sha_core/n10864_1 )
);
defparam \top/processor/sha_core/n10864_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10863_s  (
	.I0(\top/processor/sha_core/h1 [27]),
	.I1(\top/processor/sha_core/b [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10864_2 ),
	.COUT(\top/processor/sha_core/n10863_2 ),
	.SUM(\top/processor/sha_core/n10863_1 )
);
defparam \top/processor/sha_core/n10863_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10862_s  (
	.I0(\top/processor/sha_core/h1 [28]),
	.I1(\top/processor/sha_core/b [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10863_2 ),
	.COUT(\top/processor/sha_core/n10862_2 ),
	.SUM(\top/processor/sha_core/n10862_1 )
);
defparam \top/processor/sha_core/n10862_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10861_s  (
	.I0(\top/processor/sha_core/h1 [29]),
	.I1(\top/processor/sha_core/b [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10862_2 ),
	.COUT(\top/processor/sha_core/n10861_2 ),
	.SUM(\top/processor/sha_core/n10861_1 )
);
defparam \top/processor/sha_core/n10861_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10860_s  (
	.I0(\top/processor/sha_core/h1 [30]),
	.I1(\top/processor/sha_core/b [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10861_2 ),
	.COUT(\top/processor/sha_core/n10860_2 ),
	.SUM(\top/processor/sha_core/n10860_1 )
);
defparam \top/processor/sha_core/n10860_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10859_s  (
	.I0(\top/processor/sha_core/h1 [31]),
	.I1(\top/processor/sha_core/b [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10860_2 ),
	.COUT(\top/processor/sha_core/n10859_0_COUT ),
	.SUM(\top/processor/sha_core/n10859_1 )
);
defparam \top/processor/sha_core/n10859_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10923_s  (
	.I0(\top/processor/sha_core/h2 [0]),
	.I1(\top/processor/sha_core/c [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10923_2 ),
	.SUM(\top/processor/sha_core/n10923_1 )
);
defparam \top/processor/sha_core/n10923_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10922_s  (
	.I0(\top/processor/sha_core/h2 [1]),
	.I1(\top/processor/sha_core/c [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10923_2 ),
	.COUT(\top/processor/sha_core/n10922_2 ),
	.SUM(\top/processor/sha_core/n10922_1 )
);
defparam \top/processor/sha_core/n10922_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10921_s  (
	.I0(\top/processor/sha_core/h2 [2]),
	.I1(\top/processor/sha_core/c [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10922_2 ),
	.COUT(\top/processor/sha_core/n10921_2 ),
	.SUM(\top/processor/sha_core/n10921_1 )
);
defparam \top/processor/sha_core/n10921_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10920_s  (
	.I0(\top/processor/sha_core/h2 [3]),
	.I1(\top/processor/sha_core/c [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10921_2 ),
	.COUT(\top/processor/sha_core/n10920_2 ),
	.SUM(\top/processor/sha_core/n10920_1 )
);
defparam \top/processor/sha_core/n10920_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10919_s  (
	.I0(\top/processor/sha_core/h2 [4]),
	.I1(\top/processor/sha_core/c [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10920_2 ),
	.COUT(\top/processor/sha_core/n10919_2 ),
	.SUM(\top/processor/sha_core/n10919_1 )
);
defparam \top/processor/sha_core/n10919_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10918_s  (
	.I0(\top/processor/sha_core/h2 [5]),
	.I1(\top/processor/sha_core/c [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10919_2 ),
	.COUT(\top/processor/sha_core/n10918_2 ),
	.SUM(\top/processor/sha_core/n10918_1 )
);
defparam \top/processor/sha_core/n10918_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10917_s  (
	.I0(\top/processor/sha_core/h2 [6]),
	.I1(\top/processor/sha_core/c [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10918_2 ),
	.COUT(\top/processor/sha_core/n10917_2 ),
	.SUM(\top/processor/sha_core/n10917_1 )
);
defparam \top/processor/sha_core/n10917_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10916_s  (
	.I0(\top/processor/sha_core/h2 [7]),
	.I1(\top/processor/sha_core/c [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10917_2 ),
	.COUT(\top/processor/sha_core/n10916_2 ),
	.SUM(\top/processor/sha_core/n10916_1 )
);
defparam \top/processor/sha_core/n10916_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10915_s  (
	.I0(\top/processor/sha_core/h2 [8]),
	.I1(\top/processor/sha_core/c [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10916_2 ),
	.COUT(\top/processor/sha_core/n10915_2 ),
	.SUM(\top/processor/sha_core/n10915_1 )
);
defparam \top/processor/sha_core/n10915_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10914_s  (
	.I0(\top/processor/sha_core/h2 [9]),
	.I1(\top/processor/sha_core/c [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10915_2 ),
	.COUT(\top/processor/sha_core/n10914_2 ),
	.SUM(\top/processor/sha_core/n10914_1 )
);
defparam \top/processor/sha_core/n10914_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10913_s  (
	.I0(\top/processor/sha_core/h2 [10]),
	.I1(\top/processor/sha_core/c [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10914_2 ),
	.COUT(\top/processor/sha_core/n10913_2 ),
	.SUM(\top/processor/sha_core/n10913_1 )
);
defparam \top/processor/sha_core/n10913_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10912_s  (
	.I0(\top/processor/sha_core/h2 [11]),
	.I1(\top/processor/sha_core/c [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10913_2 ),
	.COUT(\top/processor/sha_core/n10912_2 ),
	.SUM(\top/processor/sha_core/n10912_1 )
);
defparam \top/processor/sha_core/n10912_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10911_s  (
	.I0(\top/processor/sha_core/h2 [12]),
	.I1(\top/processor/sha_core/c [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10912_2 ),
	.COUT(\top/processor/sha_core/n10911_2 ),
	.SUM(\top/processor/sha_core/n10911_1 )
);
defparam \top/processor/sha_core/n10911_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10910_s  (
	.I0(\top/processor/sha_core/h2 [13]),
	.I1(\top/processor/sha_core/c [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10911_2 ),
	.COUT(\top/processor/sha_core/n10910_2 ),
	.SUM(\top/processor/sha_core/n10910_1 )
);
defparam \top/processor/sha_core/n10910_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10909_s  (
	.I0(\top/processor/sha_core/h2 [14]),
	.I1(\top/processor/sha_core/c [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10910_2 ),
	.COUT(\top/processor/sha_core/n10909_2 ),
	.SUM(\top/processor/sha_core/n10909_1 )
);
defparam \top/processor/sha_core/n10909_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10908_s  (
	.I0(\top/processor/sha_core/h2 [15]),
	.I1(\top/processor/sha_core/c [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10909_2 ),
	.COUT(\top/processor/sha_core/n10908_2 ),
	.SUM(\top/processor/sha_core/n10908_1 )
);
defparam \top/processor/sha_core/n10908_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10907_s  (
	.I0(\top/processor/sha_core/h2 [16]),
	.I1(\top/processor/sha_core/c [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10908_2 ),
	.COUT(\top/processor/sha_core/n10907_2 ),
	.SUM(\top/processor/sha_core/n10907_1 )
);
defparam \top/processor/sha_core/n10907_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10906_s  (
	.I0(\top/processor/sha_core/h2 [17]),
	.I1(\top/processor/sha_core/c [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10907_2 ),
	.COUT(\top/processor/sha_core/n10906_2 ),
	.SUM(\top/processor/sha_core/n10906_1 )
);
defparam \top/processor/sha_core/n10906_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10905_s  (
	.I0(\top/processor/sha_core/h2 [18]),
	.I1(\top/processor/sha_core/c [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10906_2 ),
	.COUT(\top/processor/sha_core/n10905_2 ),
	.SUM(\top/processor/sha_core/n10905_1 )
);
defparam \top/processor/sha_core/n10905_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10904_s  (
	.I0(\top/processor/sha_core/h2 [19]),
	.I1(\top/processor/sha_core/c [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10905_2 ),
	.COUT(\top/processor/sha_core/n10904_2 ),
	.SUM(\top/processor/sha_core/n10904_1 )
);
defparam \top/processor/sha_core/n10904_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10903_s  (
	.I0(\top/processor/sha_core/h2 [20]),
	.I1(\top/processor/sha_core/c [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10904_2 ),
	.COUT(\top/processor/sha_core/n10903_2 ),
	.SUM(\top/processor/sha_core/n10903_1 )
);
defparam \top/processor/sha_core/n10903_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10902_s  (
	.I0(\top/processor/sha_core/h2 [21]),
	.I1(\top/processor/sha_core/c [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10903_2 ),
	.COUT(\top/processor/sha_core/n10902_2 ),
	.SUM(\top/processor/sha_core/n10902_1 )
);
defparam \top/processor/sha_core/n10902_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10901_s  (
	.I0(\top/processor/sha_core/h2 [22]),
	.I1(\top/processor/sha_core/c [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10902_2 ),
	.COUT(\top/processor/sha_core/n10901_2 ),
	.SUM(\top/processor/sha_core/n10901_1 )
);
defparam \top/processor/sha_core/n10901_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10900_s  (
	.I0(\top/processor/sha_core/h2 [23]),
	.I1(\top/processor/sha_core/c [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10901_2 ),
	.COUT(\top/processor/sha_core/n10900_2 ),
	.SUM(\top/processor/sha_core/n10900_1 )
);
defparam \top/processor/sha_core/n10900_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10899_s  (
	.I0(\top/processor/sha_core/h2 [24]),
	.I1(\top/processor/sha_core/c [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10900_2 ),
	.COUT(\top/processor/sha_core/n10899_2 ),
	.SUM(\top/processor/sha_core/n10899_1 )
);
defparam \top/processor/sha_core/n10899_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10898_s  (
	.I0(\top/processor/sha_core/h2 [25]),
	.I1(\top/processor/sha_core/c [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10899_2 ),
	.COUT(\top/processor/sha_core/n10898_2 ),
	.SUM(\top/processor/sha_core/n10898_1 )
);
defparam \top/processor/sha_core/n10898_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10897_s  (
	.I0(\top/processor/sha_core/h2 [26]),
	.I1(\top/processor/sha_core/c [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10898_2 ),
	.COUT(\top/processor/sha_core/n10897_2 ),
	.SUM(\top/processor/sha_core/n10897_1 )
);
defparam \top/processor/sha_core/n10897_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10896_s  (
	.I0(\top/processor/sha_core/h2 [27]),
	.I1(\top/processor/sha_core/c [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10897_2 ),
	.COUT(\top/processor/sha_core/n10896_2 ),
	.SUM(\top/processor/sha_core/n10896_1 )
);
defparam \top/processor/sha_core/n10896_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10895_s  (
	.I0(\top/processor/sha_core/h2 [28]),
	.I1(\top/processor/sha_core/c [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10896_2 ),
	.COUT(\top/processor/sha_core/n10895_2 ),
	.SUM(\top/processor/sha_core/n10895_1 )
);
defparam \top/processor/sha_core/n10895_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10894_s  (
	.I0(\top/processor/sha_core/h2 [29]),
	.I1(\top/processor/sha_core/c [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10895_2 ),
	.COUT(\top/processor/sha_core/n10894_2 ),
	.SUM(\top/processor/sha_core/n10894_1 )
);
defparam \top/processor/sha_core/n10894_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10893_s  (
	.I0(\top/processor/sha_core/h2 [30]),
	.I1(\top/processor/sha_core/c [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10894_2 ),
	.COUT(\top/processor/sha_core/n10893_2 ),
	.SUM(\top/processor/sha_core/n10893_1 )
);
defparam \top/processor/sha_core/n10893_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10892_s  (
	.I0(\top/processor/sha_core/h2 [31]),
	.I1(\top/processor/sha_core/c [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10893_2 ),
	.COUT(\top/processor/sha_core/n10892_0_COUT ),
	.SUM(\top/processor/sha_core/n10892_1 )
);
defparam \top/processor/sha_core/n10892_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10956_s  (
	.I0(\top/processor/sha_core/h3 [0]),
	.I1(\top/processor/sha_core/d [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10956_2 ),
	.SUM(\top/processor/sha_core/n10956_1 )
);
defparam \top/processor/sha_core/n10956_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10955_s  (
	.I0(\top/processor/sha_core/h3 [1]),
	.I1(\top/processor/sha_core/d [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10956_2 ),
	.COUT(\top/processor/sha_core/n10955_2 ),
	.SUM(\top/processor/sha_core/n10955_1 )
);
defparam \top/processor/sha_core/n10955_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10954_s  (
	.I0(\top/processor/sha_core/h3 [2]),
	.I1(\top/processor/sha_core/d [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10955_2 ),
	.COUT(\top/processor/sha_core/n10954_2 ),
	.SUM(\top/processor/sha_core/n10954_1 )
);
defparam \top/processor/sha_core/n10954_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10953_s  (
	.I0(\top/processor/sha_core/h3 [3]),
	.I1(\top/processor/sha_core/d [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10954_2 ),
	.COUT(\top/processor/sha_core/n10953_2 ),
	.SUM(\top/processor/sha_core/n10953_1 )
);
defparam \top/processor/sha_core/n10953_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10952_s  (
	.I0(\top/processor/sha_core/h3 [4]),
	.I1(\top/processor/sha_core/d [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10953_2 ),
	.COUT(\top/processor/sha_core/n10952_2 ),
	.SUM(\top/processor/sha_core/n10952_1 )
);
defparam \top/processor/sha_core/n10952_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10951_s  (
	.I0(\top/processor/sha_core/h3 [5]),
	.I1(\top/processor/sha_core/d [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10952_2 ),
	.COUT(\top/processor/sha_core/n10951_2 ),
	.SUM(\top/processor/sha_core/n10951_1 )
);
defparam \top/processor/sha_core/n10951_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10950_s  (
	.I0(\top/processor/sha_core/h3 [6]),
	.I1(\top/processor/sha_core/d [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10951_2 ),
	.COUT(\top/processor/sha_core/n10950_2 ),
	.SUM(\top/processor/sha_core/n10950_1 )
);
defparam \top/processor/sha_core/n10950_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10949_s  (
	.I0(\top/processor/sha_core/h3 [7]),
	.I1(\top/processor/sha_core/d [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10950_2 ),
	.COUT(\top/processor/sha_core/n10949_2 ),
	.SUM(\top/processor/sha_core/n10949_1 )
);
defparam \top/processor/sha_core/n10949_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10948_s  (
	.I0(\top/processor/sha_core/h3 [8]),
	.I1(\top/processor/sha_core/d [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10949_2 ),
	.COUT(\top/processor/sha_core/n10948_2 ),
	.SUM(\top/processor/sha_core/n10948_1 )
);
defparam \top/processor/sha_core/n10948_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10947_s  (
	.I0(\top/processor/sha_core/h3 [9]),
	.I1(\top/processor/sha_core/d [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10948_2 ),
	.COUT(\top/processor/sha_core/n10947_2 ),
	.SUM(\top/processor/sha_core/n10947_1 )
);
defparam \top/processor/sha_core/n10947_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10946_s  (
	.I0(\top/processor/sha_core/h3 [10]),
	.I1(\top/processor/sha_core/d [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10947_2 ),
	.COUT(\top/processor/sha_core/n10946_2 ),
	.SUM(\top/processor/sha_core/n10946_1 )
);
defparam \top/processor/sha_core/n10946_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10945_s  (
	.I0(\top/processor/sha_core/h3 [11]),
	.I1(\top/processor/sha_core/d [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10946_2 ),
	.COUT(\top/processor/sha_core/n10945_2 ),
	.SUM(\top/processor/sha_core/n10945_1 )
);
defparam \top/processor/sha_core/n10945_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10944_s  (
	.I0(\top/processor/sha_core/h3 [12]),
	.I1(\top/processor/sha_core/d [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10945_2 ),
	.COUT(\top/processor/sha_core/n10944_2 ),
	.SUM(\top/processor/sha_core/n10944_1 )
);
defparam \top/processor/sha_core/n10944_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10943_s  (
	.I0(\top/processor/sha_core/h3 [13]),
	.I1(\top/processor/sha_core/d [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10944_2 ),
	.COUT(\top/processor/sha_core/n10943_2 ),
	.SUM(\top/processor/sha_core/n10943_1 )
);
defparam \top/processor/sha_core/n10943_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10942_s  (
	.I0(\top/processor/sha_core/h3 [14]),
	.I1(\top/processor/sha_core/d [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10943_2 ),
	.COUT(\top/processor/sha_core/n10942_2 ),
	.SUM(\top/processor/sha_core/n10942_1 )
);
defparam \top/processor/sha_core/n10942_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10941_s  (
	.I0(\top/processor/sha_core/h3 [15]),
	.I1(\top/processor/sha_core/d [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10942_2 ),
	.COUT(\top/processor/sha_core/n10941_2 ),
	.SUM(\top/processor/sha_core/n10941_1 )
);
defparam \top/processor/sha_core/n10941_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10940_s  (
	.I0(\top/processor/sha_core/h3 [16]),
	.I1(\top/processor/sha_core/d [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10941_2 ),
	.COUT(\top/processor/sha_core/n10940_2 ),
	.SUM(\top/processor/sha_core/n10940_1 )
);
defparam \top/processor/sha_core/n10940_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10939_s  (
	.I0(\top/processor/sha_core/h3 [17]),
	.I1(\top/processor/sha_core/d [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10940_2 ),
	.COUT(\top/processor/sha_core/n10939_2 ),
	.SUM(\top/processor/sha_core/n10939_1 )
);
defparam \top/processor/sha_core/n10939_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10938_s  (
	.I0(\top/processor/sha_core/h3 [18]),
	.I1(\top/processor/sha_core/d [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10939_2 ),
	.COUT(\top/processor/sha_core/n10938_2 ),
	.SUM(\top/processor/sha_core/n10938_1 )
);
defparam \top/processor/sha_core/n10938_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10937_s  (
	.I0(\top/processor/sha_core/h3 [19]),
	.I1(\top/processor/sha_core/d [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10938_2 ),
	.COUT(\top/processor/sha_core/n10937_2 ),
	.SUM(\top/processor/sha_core/n10937_1 )
);
defparam \top/processor/sha_core/n10937_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10936_s  (
	.I0(\top/processor/sha_core/h3 [20]),
	.I1(\top/processor/sha_core/d [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10937_2 ),
	.COUT(\top/processor/sha_core/n10936_2 ),
	.SUM(\top/processor/sha_core/n10936_1 )
);
defparam \top/processor/sha_core/n10936_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10935_s  (
	.I0(\top/processor/sha_core/h3 [21]),
	.I1(\top/processor/sha_core/d [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10936_2 ),
	.COUT(\top/processor/sha_core/n10935_2 ),
	.SUM(\top/processor/sha_core/n10935_1 )
);
defparam \top/processor/sha_core/n10935_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10934_s  (
	.I0(\top/processor/sha_core/h3 [22]),
	.I1(\top/processor/sha_core/d [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10935_2 ),
	.COUT(\top/processor/sha_core/n10934_2 ),
	.SUM(\top/processor/sha_core/n10934_1 )
);
defparam \top/processor/sha_core/n10934_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10933_s  (
	.I0(\top/processor/sha_core/h3 [23]),
	.I1(\top/processor/sha_core/d [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10934_2 ),
	.COUT(\top/processor/sha_core/n10933_2 ),
	.SUM(\top/processor/sha_core/n10933_1 )
);
defparam \top/processor/sha_core/n10933_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10932_s  (
	.I0(\top/processor/sha_core/h3 [24]),
	.I1(\top/processor/sha_core/d [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10933_2 ),
	.COUT(\top/processor/sha_core/n10932_2 ),
	.SUM(\top/processor/sha_core/n10932_1 )
);
defparam \top/processor/sha_core/n10932_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10931_s  (
	.I0(\top/processor/sha_core/h3 [25]),
	.I1(\top/processor/sha_core/d [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10932_2 ),
	.COUT(\top/processor/sha_core/n10931_2 ),
	.SUM(\top/processor/sha_core/n10931_1 )
);
defparam \top/processor/sha_core/n10931_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10930_s  (
	.I0(\top/processor/sha_core/h3 [26]),
	.I1(\top/processor/sha_core/d [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10931_2 ),
	.COUT(\top/processor/sha_core/n10930_2 ),
	.SUM(\top/processor/sha_core/n10930_1 )
);
defparam \top/processor/sha_core/n10930_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10929_s  (
	.I0(\top/processor/sha_core/h3 [27]),
	.I1(\top/processor/sha_core/d [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10930_2 ),
	.COUT(\top/processor/sha_core/n10929_2 ),
	.SUM(\top/processor/sha_core/n10929_1 )
);
defparam \top/processor/sha_core/n10929_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10928_s  (
	.I0(\top/processor/sha_core/h3 [28]),
	.I1(\top/processor/sha_core/d [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10929_2 ),
	.COUT(\top/processor/sha_core/n10928_2 ),
	.SUM(\top/processor/sha_core/n10928_1 )
);
defparam \top/processor/sha_core/n10928_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10927_s  (
	.I0(\top/processor/sha_core/h3 [29]),
	.I1(\top/processor/sha_core/d [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10928_2 ),
	.COUT(\top/processor/sha_core/n10927_2 ),
	.SUM(\top/processor/sha_core/n10927_1 )
);
defparam \top/processor/sha_core/n10927_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10926_s  (
	.I0(\top/processor/sha_core/h3 [30]),
	.I1(\top/processor/sha_core/d [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10927_2 ),
	.COUT(\top/processor/sha_core/n10926_2 ),
	.SUM(\top/processor/sha_core/n10926_1 )
);
defparam \top/processor/sha_core/n10926_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10925_s  (
	.I0(\top/processor/sha_core/h3 [31]),
	.I1(\top/processor/sha_core/d [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10926_2 ),
	.COUT(\top/processor/sha_core/n10925_0_COUT ),
	.SUM(\top/processor/sha_core/n10925_1 )
);
defparam \top/processor/sha_core/n10925_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10989_s  (
	.I0(\top/processor/sha_core/h4 [0]),
	.I1(\top/processor/sha_core/e [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10989_2 ),
	.SUM(\top/processor/sha_core/n10989_1 )
);
defparam \top/processor/sha_core/n10989_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10988_s  (
	.I0(\top/processor/sha_core/h4 [1]),
	.I1(\top/processor/sha_core/e [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10989_2 ),
	.COUT(\top/processor/sha_core/n10988_2 ),
	.SUM(\top/processor/sha_core/n10988_1 )
);
defparam \top/processor/sha_core/n10988_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10987_s  (
	.I0(\top/processor/sha_core/h4 [2]),
	.I1(\top/processor/sha_core/e [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10988_2 ),
	.COUT(\top/processor/sha_core/n10987_2 ),
	.SUM(\top/processor/sha_core/n10987_1 )
);
defparam \top/processor/sha_core/n10987_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10986_s  (
	.I0(\top/processor/sha_core/h4 [3]),
	.I1(\top/processor/sha_core/e [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10987_2 ),
	.COUT(\top/processor/sha_core/n10986_2 ),
	.SUM(\top/processor/sha_core/n10986_1 )
);
defparam \top/processor/sha_core/n10986_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10985_s  (
	.I0(\top/processor/sha_core/h4 [4]),
	.I1(\top/processor/sha_core/e [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10986_2 ),
	.COUT(\top/processor/sha_core/n10985_2 ),
	.SUM(\top/processor/sha_core/n10985_1 )
);
defparam \top/processor/sha_core/n10985_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10984_s  (
	.I0(\top/processor/sha_core/h4 [5]),
	.I1(\top/processor/sha_core/e [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10985_2 ),
	.COUT(\top/processor/sha_core/n10984_2 ),
	.SUM(\top/processor/sha_core/n10984_1 )
);
defparam \top/processor/sha_core/n10984_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10983_s  (
	.I0(\top/processor/sha_core/h4 [6]),
	.I1(\top/processor/sha_core/e [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10984_2 ),
	.COUT(\top/processor/sha_core/n10983_2 ),
	.SUM(\top/processor/sha_core/n10983_1 )
);
defparam \top/processor/sha_core/n10983_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10982_s  (
	.I0(\top/processor/sha_core/h4 [7]),
	.I1(\top/processor/sha_core/e [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10983_2 ),
	.COUT(\top/processor/sha_core/n10982_2 ),
	.SUM(\top/processor/sha_core/n10982_1 )
);
defparam \top/processor/sha_core/n10982_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10981_s  (
	.I0(\top/processor/sha_core/h4 [8]),
	.I1(\top/processor/sha_core/e [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10982_2 ),
	.COUT(\top/processor/sha_core/n10981_2 ),
	.SUM(\top/processor/sha_core/n10981_1 )
);
defparam \top/processor/sha_core/n10981_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10980_s  (
	.I0(\top/processor/sha_core/h4 [9]),
	.I1(\top/processor/sha_core/e [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10981_2 ),
	.COUT(\top/processor/sha_core/n10980_2 ),
	.SUM(\top/processor/sha_core/n10980_1 )
);
defparam \top/processor/sha_core/n10980_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10979_s  (
	.I0(\top/processor/sha_core/h4 [10]),
	.I1(\top/processor/sha_core/e [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10980_2 ),
	.COUT(\top/processor/sha_core/n10979_2 ),
	.SUM(\top/processor/sha_core/n10979_1 )
);
defparam \top/processor/sha_core/n10979_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10978_s  (
	.I0(\top/processor/sha_core/h4 [11]),
	.I1(\top/processor/sha_core/e [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10979_2 ),
	.COUT(\top/processor/sha_core/n10978_2 ),
	.SUM(\top/processor/sha_core/n10978_1 )
);
defparam \top/processor/sha_core/n10978_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10977_s  (
	.I0(\top/processor/sha_core/h4 [12]),
	.I1(\top/processor/sha_core/e [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10978_2 ),
	.COUT(\top/processor/sha_core/n10977_2 ),
	.SUM(\top/processor/sha_core/n10977_1 )
);
defparam \top/processor/sha_core/n10977_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10976_s  (
	.I0(\top/processor/sha_core/h4 [13]),
	.I1(\top/processor/sha_core/e [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10977_2 ),
	.COUT(\top/processor/sha_core/n10976_2 ),
	.SUM(\top/processor/sha_core/n10976_1 )
);
defparam \top/processor/sha_core/n10976_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10975_s  (
	.I0(\top/processor/sha_core/h4 [14]),
	.I1(\top/processor/sha_core/e [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10976_2 ),
	.COUT(\top/processor/sha_core/n10975_2 ),
	.SUM(\top/processor/sha_core/n10975_1 )
);
defparam \top/processor/sha_core/n10975_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10974_s  (
	.I0(\top/processor/sha_core/h4 [15]),
	.I1(\top/processor/sha_core/e [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10975_2 ),
	.COUT(\top/processor/sha_core/n10974_2 ),
	.SUM(\top/processor/sha_core/n10974_1 )
);
defparam \top/processor/sha_core/n10974_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10973_s  (
	.I0(\top/processor/sha_core/h4 [16]),
	.I1(\top/processor/sha_core/e [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10974_2 ),
	.COUT(\top/processor/sha_core/n10973_2 ),
	.SUM(\top/processor/sha_core/n10973_1 )
);
defparam \top/processor/sha_core/n10973_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10972_s  (
	.I0(\top/processor/sha_core/h4 [17]),
	.I1(\top/processor/sha_core/e [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10973_2 ),
	.COUT(\top/processor/sha_core/n10972_2 ),
	.SUM(\top/processor/sha_core/n10972_1 )
);
defparam \top/processor/sha_core/n10972_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10971_s  (
	.I0(\top/processor/sha_core/h4 [18]),
	.I1(\top/processor/sha_core/e [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10972_2 ),
	.COUT(\top/processor/sha_core/n10971_2 ),
	.SUM(\top/processor/sha_core/n10971_1 )
);
defparam \top/processor/sha_core/n10971_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10970_s  (
	.I0(\top/processor/sha_core/h4 [19]),
	.I1(\top/processor/sha_core/e [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10971_2 ),
	.COUT(\top/processor/sha_core/n10970_2 ),
	.SUM(\top/processor/sha_core/n10970_1 )
);
defparam \top/processor/sha_core/n10970_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10969_s  (
	.I0(\top/processor/sha_core/h4 [20]),
	.I1(\top/processor/sha_core/e [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10970_2 ),
	.COUT(\top/processor/sha_core/n10969_2 ),
	.SUM(\top/processor/sha_core/n10969_1 )
);
defparam \top/processor/sha_core/n10969_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10968_s  (
	.I0(\top/processor/sha_core/h4 [21]),
	.I1(\top/processor/sha_core/e [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10969_2 ),
	.COUT(\top/processor/sha_core/n10968_2 ),
	.SUM(\top/processor/sha_core/n10968_1 )
);
defparam \top/processor/sha_core/n10968_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10967_s  (
	.I0(\top/processor/sha_core/h4 [22]),
	.I1(\top/processor/sha_core/e [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10968_2 ),
	.COUT(\top/processor/sha_core/n10967_2 ),
	.SUM(\top/processor/sha_core/n10967_1 )
);
defparam \top/processor/sha_core/n10967_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10966_s  (
	.I0(\top/processor/sha_core/h4 [23]),
	.I1(\top/processor/sha_core/e [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10967_2 ),
	.COUT(\top/processor/sha_core/n10966_2 ),
	.SUM(\top/processor/sha_core/n10966_1 )
);
defparam \top/processor/sha_core/n10966_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10965_s  (
	.I0(\top/processor/sha_core/h4 [24]),
	.I1(\top/processor/sha_core/e [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10966_2 ),
	.COUT(\top/processor/sha_core/n10965_2 ),
	.SUM(\top/processor/sha_core/n10965_1 )
);
defparam \top/processor/sha_core/n10965_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10964_s  (
	.I0(\top/processor/sha_core/h4 [25]),
	.I1(\top/processor/sha_core/e [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10965_2 ),
	.COUT(\top/processor/sha_core/n10964_2 ),
	.SUM(\top/processor/sha_core/n10964_1 )
);
defparam \top/processor/sha_core/n10964_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10963_s  (
	.I0(\top/processor/sha_core/h4 [26]),
	.I1(\top/processor/sha_core/e [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10964_2 ),
	.COUT(\top/processor/sha_core/n10963_2 ),
	.SUM(\top/processor/sha_core/n10963_1 )
);
defparam \top/processor/sha_core/n10963_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10962_s  (
	.I0(\top/processor/sha_core/h4 [27]),
	.I1(\top/processor/sha_core/e [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10963_2 ),
	.COUT(\top/processor/sha_core/n10962_2 ),
	.SUM(\top/processor/sha_core/n10962_1 )
);
defparam \top/processor/sha_core/n10962_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10961_s  (
	.I0(\top/processor/sha_core/h4 [28]),
	.I1(\top/processor/sha_core/e [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10962_2 ),
	.COUT(\top/processor/sha_core/n10961_2 ),
	.SUM(\top/processor/sha_core/n10961_1 )
);
defparam \top/processor/sha_core/n10961_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10960_s  (
	.I0(\top/processor/sha_core/h4 [29]),
	.I1(\top/processor/sha_core/e [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10961_2 ),
	.COUT(\top/processor/sha_core/n10960_2 ),
	.SUM(\top/processor/sha_core/n10960_1 )
);
defparam \top/processor/sha_core/n10960_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10959_s  (
	.I0(\top/processor/sha_core/h4 [30]),
	.I1(\top/processor/sha_core/e [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10960_2 ),
	.COUT(\top/processor/sha_core/n10959_2 ),
	.SUM(\top/processor/sha_core/n10959_1 )
);
defparam \top/processor/sha_core/n10959_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10958_s  (
	.I0(\top/processor/sha_core/h4 [31]),
	.I1(\top/processor/sha_core/e [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10959_2 ),
	.COUT(\top/processor/sha_core/n10958_0_COUT ),
	.SUM(\top/processor/sha_core/n10958_1 )
);
defparam \top/processor/sha_core/n10958_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11022_s  (
	.I0(\top/processor/sha_core/h5 [0]),
	.I1(\top/processor/sha_core/f [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n11022_2 ),
	.SUM(\top/processor/sha_core/n11022_1 )
);
defparam \top/processor/sha_core/n11022_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11021_s  (
	.I0(\top/processor/sha_core/h5 [1]),
	.I1(\top/processor/sha_core/f [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11022_2 ),
	.COUT(\top/processor/sha_core/n11021_2 ),
	.SUM(\top/processor/sha_core/n11021_1 )
);
defparam \top/processor/sha_core/n11021_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11020_s  (
	.I0(\top/processor/sha_core/h5 [2]),
	.I1(\top/processor/sha_core/f [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11021_2 ),
	.COUT(\top/processor/sha_core/n11020_2 ),
	.SUM(\top/processor/sha_core/n11020_1 )
);
defparam \top/processor/sha_core/n11020_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11019_s  (
	.I0(\top/processor/sha_core/h5 [3]),
	.I1(\top/processor/sha_core/f [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11020_2 ),
	.COUT(\top/processor/sha_core/n11019_2 ),
	.SUM(\top/processor/sha_core/n11019_1 )
);
defparam \top/processor/sha_core/n11019_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11018_s  (
	.I0(\top/processor/sha_core/h5 [4]),
	.I1(\top/processor/sha_core/f [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11019_2 ),
	.COUT(\top/processor/sha_core/n11018_2 ),
	.SUM(\top/processor/sha_core/n11018_1 )
);
defparam \top/processor/sha_core/n11018_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11017_s  (
	.I0(\top/processor/sha_core/h5 [5]),
	.I1(\top/processor/sha_core/f [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11018_2 ),
	.COUT(\top/processor/sha_core/n11017_2 ),
	.SUM(\top/processor/sha_core/n11017_1 )
);
defparam \top/processor/sha_core/n11017_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11016_s  (
	.I0(\top/processor/sha_core/h5 [6]),
	.I1(\top/processor/sha_core/f [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11017_2 ),
	.COUT(\top/processor/sha_core/n11016_2 ),
	.SUM(\top/processor/sha_core/n11016_1 )
);
defparam \top/processor/sha_core/n11016_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11015_s  (
	.I0(\top/processor/sha_core/h5 [7]),
	.I1(\top/processor/sha_core/f [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11016_2 ),
	.COUT(\top/processor/sha_core/n11015_2 ),
	.SUM(\top/processor/sha_core/n11015_1 )
);
defparam \top/processor/sha_core/n11015_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11014_s  (
	.I0(\top/processor/sha_core/h5 [8]),
	.I1(\top/processor/sha_core/f [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11015_2 ),
	.COUT(\top/processor/sha_core/n11014_2 ),
	.SUM(\top/processor/sha_core/n11014_1 )
);
defparam \top/processor/sha_core/n11014_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11013_s  (
	.I0(\top/processor/sha_core/h5 [9]),
	.I1(\top/processor/sha_core/f [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11014_2 ),
	.COUT(\top/processor/sha_core/n11013_2 ),
	.SUM(\top/processor/sha_core/n11013_1 )
);
defparam \top/processor/sha_core/n11013_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11012_s  (
	.I0(\top/processor/sha_core/h5 [10]),
	.I1(\top/processor/sha_core/f [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11013_2 ),
	.COUT(\top/processor/sha_core/n11012_2 ),
	.SUM(\top/processor/sha_core/n11012_1 )
);
defparam \top/processor/sha_core/n11012_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11011_s  (
	.I0(\top/processor/sha_core/h5 [11]),
	.I1(\top/processor/sha_core/f [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11012_2 ),
	.COUT(\top/processor/sha_core/n11011_2 ),
	.SUM(\top/processor/sha_core/n11011_1 )
);
defparam \top/processor/sha_core/n11011_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11010_s  (
	.I0(\top/processor/sha_core/h5 [12]),
	.I1(\top/processor/sha_core/f [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11011_2 ),
	.COUT(\top/processor/sha_core/n11010_2 ),
	.SUM(\top/processor/sha_core/n11010_1 )
);
defparam \top/processor/sha_core/n11010_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11009_s  (
	.I0(\top/processor/sha_core/h5 [13]),
	.I1(\top/processor/sha_core/f [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11010_2 ),
	.COUT(\top/processor/sha_core/n11009_2 ),
	.SUM(\top/processor/sha_core/n11009_1 )
);
defparam \top/processor/sha_core/n11009_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11008_s  (
	.I0(\top/processor/sha_core/h5 [14]),
	.I1(\top/processor/sha_core/f [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11009_2 ),
	.COUT(\top/processor/sha_core/n11008_2 ),
	.SUM(\top/processor/sha_core/n11008_1 )
);
defparam \top/processor/sha_core/n11008_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11007_s  (
	.I0(\top/processor/sha_core/h5 [15]),
	.I1(\top/processor/sha_core/f [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11008_2 ),
	.COUT(\top/processor/sha_core/n11007_2 ),
	.SUM(\top/processor/sha_core/n11007_1 )
);
defparam \top/processor/sha_core/n11007_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11006_s  (
	.I0(\top/processor/sha_core/h5 [16]),
	.I1(\top/processor/sha_core/f [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11007_2 ),
	.COUT(\top/processor/sha_core/n11006_2 ),
	.SUM(\top/processor/sha_core/n11006_1 )
);
defparam \top/processor/sha_core/n11006_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11005_s  (
	.I0(\top/processor/sha_core/h5 [17]),
	.I1(\top/processor/sha_core/f [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11006_2 ),
	.COUT(\top/processor/sha_core/n11005_2 ),
	.SUM(\top/processor/sha_core/n11005_1 )
);
defparam \top/processor/sha_core/n11005_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11004_s  (
	.I0(\top/processor/sha_core/h5 [18]),
	.I1(\top/processor/sha_core/f [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11005_2 ),
	.COUT(\top/processor/sha_core/n11004_2 ),
	.SUM(\top/processor/sha_core/n11004_1 )
);
defparam \top/processor/sha_core/n11004_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11003_s  (
	.I0(\top/processor/sha_core/h5 [19]),
	.I1(\top/processor/sha_core/f [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11004_2 ),
	.COUT(\top/processor/sha_core/n11003_2 ),
	.SUM(\top/processor/sha_core/n11003_1 )
);
defparam \top/processor/sha_core/n11003_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11002_s  (
	.I0(\top/processor/sha_core/h5 [20]),
	.I1(\top/processor/sha_core/f [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11003_2 ),
	.COUT(\top/processor/sha_core/n11002_2 ),
	.SUM(\top/processor/sha_core/n11002_1 )
);
defparam \top/processor/sha_core/n11002_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11001_s  (
	.I0(\top/processor/sha_core/h5 [21]),
	.I1(\top/processor/sha_core/f [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11002_2 ),
	.COUT(\top/processor/sha_core/n11001_2 ),
	.SUM(\top/processor/sha_core/n11001_1 )
);
defparam \top/processor/sha_core/n11001_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11000_s  (
	.I0(\top/processor/sha_core/h5 [22]),
	.I1(\top/processor/sha_core/f [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11001_2 ),
	.COUT(\top/processor/sha_core/n11000_2 ),
	.SUM(\top/processor/sha_core/n11000_1 )
);
defparam \top/processor/sha_core/n11000_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10999_s  (
	.I0(\top/processor/sha_core/h5 [23]),
	.I1(\top/processor/sha_core/f [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11000_2 ),
	.COUT(\top/processor/sha_core/n10999_2 ),
	.SUM(\top/processor/sha_core/n10999_1 )
);
defparam \top/processor/sha_core/n10999_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10998_s  (
	.I0(\top/processor/sha_core/h5 [24]),
	.I1(\top/processor/sha_core/f [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10999_2 ),
	.COUT(\top/processor/sha_core/n10998_2 ),
	.SUM(\top/processor/sha_core/n10998_1 )
);
defparam \top/processor/sha_core/n10998_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10997_s  (
	.I0(\top/processor/sha_core/h5 [25]),
	.I1(\top/processor/sha_core/f [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10998_2 ),
	.COUT(\top/processor/sha_core/n10997_2 ),
	.SUM(\top/processor/sha_core/n10997_1 )
);
defparam \top/processor/sha_core/n10997_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10996_s  (
	.I0(\top/processor/sha_core/h5 [26]),
	.I1(\top/processor/sha_core/f [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10997_2 ),
	.COUT(\top/processor/sha_core/n10996_2 ),
	.SUM(\top/processor/sha_core/n10996_1 )
);
defparam \top/processor/sha_core/n10996_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10995_s  (
	.I0(\top/processor/sha_core/h5 [27]),
	.I1(\top/processor/sha_core/f [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10996_2 ),
	.COUT(\top/processor/sha_core/n10995_2 ),
	.SUM(\top/processor/sha_core/n10995_1 )
);
defparam \top/processor/sha_core/n10995_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10994_s  (
	.I0(\top/processor/sha_core/h5 [28]),
	.I1(\top/processor/sha_core/f [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10995_2 ),
	.COUT(\top/processor/sha_core/n10994_2 ),
	.SUM(\top/processor/sha_core/n10994_1 )
);
defparam \top/processor/sha_core/n10994_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10993_s  (
	.I0(\top/processor/sha_core/h5 [29]),
	.I1(\top/processor/sha_core/f [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10994_2 ),
	.COUT(\top/processor/sha_core/n10993_2 ),
	.SUM(\top/processor/sha_core/n10993_1 )
);
defparam \top/processor/sha_core/n10993_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10992_s  (
	.I0(\top/processor/sha_core/h5 [30]),
	.I1(\top/processor/sha_core/f [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10993_2 ),
	.COUT(\top/processor/sha_core/n10992_2 ),
	.SUM(\top/processor/sha_core/n10992_1 )
);
defparam \top/processor/sha_core/n10992_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10991_s  (
	.I0(\top/processor/sha_core/h5 [31]),
	.I1(\top/processor/sha_core/f [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10992_2 ),
	.COUT(\top/processor/sha_core/n10991_0_COUT ),
	.SUM(\top/processor/sha_core/n10991_1 )
);
defparam \top/processor/sha_core/n10991_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11055_s  (
	.I0(\top/processor/sha_core/h6 [0]),
	.I1(\top/processor/sha_core/g [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n11055_2 ),
	.SUM(\top/processor/sha_core/n11055_1 )
);
defparam \top/processor/sha_core/n11055_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11054_s  (
	.I0(\top/processor/sha_core/h6 [1]),
	.I1(\top/processor/sha_core/g [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11055_2 ),
	.COUT(\top/processor/sha_core/n11054_2 ),
	.SUM(\top/processor/sha_core/n11054_1 )
);
defparam \top/processor/sha_core/n11054_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11053_s  (
	.I0(\top/processor/sha_core/h6 [2]),
	.I1(\top/processor/sha_core/g [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11054_2 ),
	.COUT(\top/processor/sha_core/n11053_2 ),
	.SUM(\top/processor/sha_core/n11053_1 )
);
defparam \top/processor/sha_core/n11053_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11052_s  (
	.I0(\top/processor/sha_core/h6 [3]),
	.I1(\top/processor/sha_core/g [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11053_2 ),
	.COUT(\top/processor/sha_core/n11052_2 ),
	.SUM(\top/processor/sha_core/n11052_1 )
);
defparam \top/processor/sha_core/n11052_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11051_s  (
	.I0(\top/processor/sha_core/h6 [4]),
	.I1(\top/processor/sha_core/g [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11052_2 ),
	.COUT(\top/processor/sha_core/n11051_2 ),
	.SUM(\top/processor/sha_core/n11051_1 )
);
defparam \top/processor/sha_core/n11051_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11050_s  (
	.I0(\top/processor/sha_core/h6 [5]),
	.I1(\top/processor/sha_core/g [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11051_2 ),
	.COUT(\top/processor/sha_core/n11050_2 ),
	.SUM(\top/processor/sha_core/n11050_1 )
);
defparam \top/processor/sha_core/n11050_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11049_s  (
	.I0(\top/processor/sha_core/h6 [6]),
	.I1(\top/processor/sha_core/g [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11050_2 ),
	.COUT(\top/processor/sha_core/n11049_2 ),
	.SUM(\top/processor/sha_core/n11049_1 )
);
defparam \top/processor/sha_core/n11049_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11048_s  (
	.I0(\top/processor/sha_core/h6 [7]),
	.I1(\top/processor/sha_core/g [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11049_2 ),
	.COUT(\top/processor/sha_core/n11048_2 ),
	.SUM(\top/processor/sha_core/n11048_1 )
);
defparam \top/processor/sha_core/n11048_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11047_s  (
	.I0(\top/processor/sha_core/h6 [8]),
	.I1(\top/processor/sha_core/g [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11048_2 ),
	.COUT(\top/processor/sha_core/n11047_2 ),
	.SUM(\top/processor/sha_core/n11047_1 )
);
defparam \top/processor/sha_core/n11047_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11046_s  (
	.I0(\top/processor/sha_core/h6 [9]),
	.I1(\top/processor/sha_core/g [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11047_2 ),
	.COUT(\top/processor/sha_core/n11046_2 ),
	.SUM(\top/processor/sha_core/n11046_1 )
);
defparam \top/processor/sha_core/n11046_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11045_s  (
	.I0(\top/processor/sha_core/h6 [10]),
	.I1(\top/processor/sha_core/g [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11046_2 ),
	.COUT(\top/processor/sha_core/n11045_2 ),
	.SUM(\top/processor/sha_core/n11045_1 )
);
defparam \top/processor/sha_core/n11045_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11044_s  (
	.I0(\top/processor/sha_core/h6 [11]),
	.I1(\top/processor/sha_core/g [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11045_2 ),
	.COUT(\top/processor/sha_core/n11044_2 ),
	.SUM(\top/processor/sha_core/n11044_1 )
);
defparam \top/processor/sha_core/n11044_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11043_s  (
	.I0(\top/processor/sha_core/h6 [12]),
	.I1(\top/processor/sha_core/g [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11044_2 ),
	.COUT(\top/processor/sha_core/n11043_2 ),
	.SUM(\top/processor/sha_core/n11043_1 )
);
defparam \top/processor/sha_core/n11043_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11042_s  (
	.I0(\top/processor/sha_core/h6 [13]),
	.I1(\top/processor/sha_core/g [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11043_2 ),
	.COUT(\top/processor/sha_core/n11042_2 ),
	.SUM(\top/processor/sha_core/n11042_1 )
);
defparam \top/processor/sha_core/n11042_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11041_s  (
	.I0(\top/processor/sha_core/h6 [14]),
	.I1(\top/processor/sha_core/g [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11042_2 ),
	.COUT(\top/processor/sha_core/n11041_2 ),
	.SUM(\top/processor/sha_core/n11041_1 )
);
defparam \top/processor/sha_core/n11041_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11040_s  (
	.I0(\top/processor/sha_core/h6 [15]),
	.I1(\top/processor/sha_core/g [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11041_2 ),
	.COUT(\top/processor/sha_core/n11040_2 ),
	.SUM(\top/processor/sha_core/n11040_1 )
);
defparam \top/processor/sha_core/n11040_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11039_s  (
	.I0(\top/processor/sha_core/h6 [16]),
	.I1(\top/processor/sha_core/g [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11040_2 ),
	.COUT(\top/processor/sha_core/n11039_2 ),
	.SUM(\top/processor/sha_core/n11039_1 )
);
defparam \top/processor/sha_core/n11039_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11038_s  (
	.I0(\top/processor/sha_core/h6 [17]),
	.I1(\top/processor/sha_core/g [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11039_2 ),
	.COUT(\top/processor/sha_core/n11038_2 ),
	.SUM(\top/processor/sha_core/n11038_1 )
);
defparam \top/processor/sha_core/n11038_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11037_s  (
	.I0(\top/processor/sha_core/h6 [18]),
	.I1(\top/processor/sha_core/g [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11038_2 ),
	.COUT(\top/processor/sha_core/n11037_2 ),
	.SUM(\top/processor/sha_core/n11037_1 )
);
defparam \top/processor/sha_core/n11037_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11036_s  (
	.I0(\top/processor/sha_core/h6 [19]),
	.I1(\top/processor/sha_core/g [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11037_2 ),
	.COUT(\top/processor/sha_core/n11036_2 ),
	.SUM(\top/processor/sha_core/n11036_1 )
);
defparam \top/processor/sha_core/n11036_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11035_s  (
	.I0(\top/processor/sha_core/h6 [20]),
	.I1(\top/processor/sha_core/g [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11036_2 ),
	.COUT(\top/processor/sha_core/n11035_2 ),
	.SUM(\top/processor/sha_core/n11035_1 )
);
defparam \top/processor/sha_core/n11035_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11034_s  (
	.I0(\top/processor/sha_core/h6 [21]),
	.I1(\top/processor/sha_core/g [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11035_2 ),
	.COUT(\top/processor/sha_core/n11034_2 ),
	.SUM(\top/processor/sha_core/n11034_1 )
);
defparam \top/processor/sha_core/n11034_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11033_s  (
	.I0(\top/processor/sha_core/h6 [22]),
	.I1(\top/processor/sha_core/g [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11034_2 ),
	.COUT(\top/processor/sha_core/n11033_2 ),
	.SUM(\top/processor/sha_core/n11033_1 )
);
defparam \top/processor/sha_core/n11033_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11032_s  (
	.I0(\top/processor/sha_core/h6 [23]),
	.I1(\top/processor/sha_core/g [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11033_2 ),
	.COUT(\top/processor/sha_core/n11032_2 ),
	.SUM(\top/processor/sha_core/n11032_1 )
);
defparam \top/processor/sha_core/n11032_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11031_s  (
	.I0(\top/processor/sha_core/h6 [24]),
	.I1(\top/processor/sha_core/g [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11032_2 ),
	.COUT(\top/processor/sha_core/n11031_2 ),
	.SUM(\top/processor/sha_core/n11031_1 )
);
defparam \top/processor/sha_core/n11031_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11030_s  (
	.I0(\top/processor/sha_core/h6 [25]),
	.I1(\top/processor/sha_core/g [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11031_2 ),
	.COUT(\top/processor/sha_core/n11030_2 ),
	.SUM(\top/processor/sha_core/n11030_1 )
);
defparam \top/processor/sha_core/n11030_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11029_s  (
	.I0(\top/processor/sha_core/h6 [26]),
	.I1(\top/processor/sha_core/g [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11030_2 ),
	.COUT(\top/processor/sha_core/n11029_2 ),
	.SUM(\top/processor/sha_core/n11029_1 )
);
defparam \top/processor/sha_core/n11029_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11028_s  (
	.I0(\top/processor/sha_core/h6 [27]),
	.I1(\top/processor/sha_core/g [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11029_2 ),
	.COUT(\top/processor/sha_core/n11028_2 ),
	.SUM(\top/processor/sha_core/n11028_1 )
);
defparam \top/processor/sha_core/n11028_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11027_s  (
	.I0(\top/processor/sha_core/h6 [28]),
	.I1(\top/processor/sha_core/g [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11028_2 ),
	.COUT(\top/processor/sha_core/n11027_2 ),
	.SUM(\top/processor/sha_core/n11027_1 )
);
defparam \top/processor/sha_core/n11027_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11026_s  (
	.I0(\top/processor/sha_core/h6 [29]),
	.I1(\top/processor/sha_core/g [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11027_2 ),
	.COUT(\top/processor/sha_core/n11026_2 ),
	.SUM(\top/processor/sha_core/n11026_1 )
);
defparam \top/processor/sha_core/n11026_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11025_s  (
	.I0(\top/processor/sha_core/h6 [30]),
	.I1(\top/processor/sha_core/g [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11026_2 ),
	.COUT(\top/processor/sha_core/n11025_2 ),
	.SUM(\top/processor/sha_core/n11025_1 )
);
defparam \top/processor/sha_core/n11025_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11024_s  (
	.I0(\top/processor/sha_core/h6 [31]),
	.I1(\top/processor/sha_core/g [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11025_2 ),
	.COUT(\top/processor/sha_core/n11024_0_COUT ),
	.SUM(\top/processor/sha_core/n11024_1 )
);
defparam \top/processor/sha_core/n11024_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11088_s  (
	.I0(\top/processor/sha_core/h7 [0]),
	.I1(\top/processor/sha_core/h [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n11088_2 ),
	.SUM(\top/processor/sha_core/n11088_1 )
);
defparam \top/processor/sha_core/n11088_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11087_s  (
	.I0(\top/processor/sha_core/h7 [1]),
	.I1(\top/processor/sha_core/h [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11088_2 ),
	.COUT(\top/processor/sha_core/n11087_2 ),
	.SUM(\top/processor/sha_core/n11087_1 )
);
defparam \top/processor/sha_core/n11087_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11086_s  (
	.I0(\top/processor/sha_core/h7 [2]),
	.I1(\top/processor/sha_core/h [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11087_2 ),
	.COUT(\top/processor/sha_core/n11086_2 ),
	.SUM(\top/processor/sha_core/n11086_1 )
);
defparam \top/processor/sha_core/n11086_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11085_s  (
	.I0(\top/processor/sha_core/h7 [3]),
	.I1(\top/processor/sha_core/h [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11086_2 ),
	.COUT(\top/processor/sha_core/n11085_2 ),
	.SUM(\top/processor/sha_core/n11085_1 )
);
defparam \top/processor/sha_core/n11085_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11084_s  (
	.I0(\top/processor/sha_core/h7 [4]),
	.I1(\top/processor/sha_core/h [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11085_2 ),
	.COUT(\top/processor/sha_core/n11084_2 ),
	.SUM(\top/processor/sha_core/n11084_1 )
);
defparam \top/processor/sha_core/n11084_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11083_s  (
	.I0(\top/processor/sha_core/h7 [5]),
	.I1(\top/processor/sha_core/h [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11084_2 ),
	.COUT(\top/processor/sha_core/n11083_2 ),
	.SUM(\top/processor/sha_core/n11083_1 )
);
defparam \top/processor/sha_core/n11083_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11082_s  (
	.I0(\top/processor/sha_core/h7 [6]),
	.I1(\top/processor/sha_core/h [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11083_2 ),
	.COUT(\top/processor/sha_core/n11082_2 ),
	.SUM(\top/processor/sha_core/n11082_1 )
);
defparam \top/processor/sha_core/n11082_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11081_s  (
	.I0(\top/processor/sha_core/h7 [7]),
	.I1(\top/processor/sha_core/h [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11082_2 ),
	.COUT(\top/processor/sha_core/n11081_2 ),
	.SUM(\top/processor/sha_core/n11081_1 )
);
defparam \top/processor/sha_core/n11081_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11080_s  (
	.I0(\top/processor/sha_core/h7 [8]),
	.I1(\top/processor/sha_core/h [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11081_2 ),
	.COUT(\top/processor/sha_core/n11080_2 ),
	.SUM(\top/processor/sha_core/n11080_1 )
);
defparam \top/processor/sha_core/n11080_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11079_s  (
	.I0(\top/processor/sha_core/h7 [9]),
	.I1(\top/processor/sha_core/h [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11080_2 ),
	.COUT(\top/processor/sha_core/n11079_2 ),
	.SUM(\top/processor/sha_core/n11079_1 )
);
defparam \top/processor/sha_core/n11079_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11078_s  (
	.I0(\top/processor/sha_core/h7 [10]),
	.I1(\top/processor/sha_core/h [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11079_2 ),
	.COUT(\top/processor/sha_core/n11078_2 ),
	.SUM(\top/processor/sha_core/n11078_1 )
);
defparam \top/processor/sha_core/n11078_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11077_s  (
	.I0(\top/processor/sha_core/h7 [11]),
	.I1(\top/processor/sha_core/h [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11078_2 ),
	.COUT(\top/processor/sha_core/n11077_2 ),
	.SUM(\top/processor/sha_core/n11077_1 )
);
defparam \top/processor/sha_core/n11077_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11076_s  (
	.I0(\top/processor/sha_core/h7 [12]),
	.I1(\top/processor/sha_core/h [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11077_2 ),
	.COUT(\top/processor/sha_core/n11076_2 ),
	.SUM(\top/processor/sha_core/n11076_1 )
);
defparam \top/processor/sha_core/n11076_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11075_s  (
	.I0(\top/processor/sha_core/h7 [13]),
	.I1(\top/processor/sha_core/h [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11076_2 ),
	.COUT(\top/processor/sha_core/n11075_2 ),
	.SUM(\top/processor/sha_core/n11075_1 )
);
defparam \top/processor/sha_core/n11075_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11074_s  (
	.I0(\top/processor/sha_core/h7 [14]),
	.I1(\top/processor/sha_core/h [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11075_2 ),
	.COUT(\top/processor/sha_core/n11074_2 ),
	.SUM(\top/processor/sha_core/n11074_1 )
);
defparam \top/processor/sha_core/n11074_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11073_s  (
	.I0(\top/processor/sha_core/h7 [15]),
	.I1(\top/processor/sha_core/h [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11074_2 ),
	.COUT(\top/processor/sha_core/n11073_2 ),
	.SUM(\top/processor/sha_core/n11073_1 )
);
defparam \top/processor/sha_core/n11073_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11072_s  (
	.I0(\top/processor/sha_core/h7 [16]),
	.I1(\top/processor/sha_core/h [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11073_2 ),
	.COUT(\top/processor/sha_core/n11072_2 ),
	.SUM(\top/processor/sha_core/n11072_1 )
);
defparam \top/processor/sha_core/n11072_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11071_s  (
	.I0(\top/processor/sha_core/h7 [17]),
	.I1(\top/processor/sha_core/h [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11072_2 ),
	.COUT(\top/processor/sha_core/n11071_2 ),
	.SUM(\top/processor/sha_core/n11071_1 )
);
defparam \top/processor/sha_core/n11071_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11070_s  (
	.I0(\top/processor/sha_core/h7 [18]),
	.I1(\top/processor/sha_core/h [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11071_2 ),
	.COUT(\top/processor/sha_core/n11070_2 ),
	.SUM(\top/processor/sha_core/n11070_1 )
);
defparam \top/processor/sha_core/n11070_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11069_s  (
	.I0(\top/processor/sha_core/h7 [19]),
	.I1(\top/processor/sha_core/h [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11070_2 ),
	.COUT(\top/processor/sha_core/n11069_2 ),
	.SUM(\top/processor/sha_core/n11069_1 )
);
defparam \top/processor/sha_core/n11069_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11068_s  (
	.I0(\top/processor/sha_core/h7 [20]),
	.I1(\top/processor/sha_core/h [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11069_2 ),
	.COUT(\top/processor/sha_core/n11068_2 ),
	.SUM(\top/processor/sha_core/n11068_1 )
);
defparam \top/processor/sha_core/n11068_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11067_s  (
	.I0(\top/processor/sha_core/h7 [21]),
	.I1(\top/processor/sha_core/h [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11068_2 ),
	.COUT(\top/processor/sha_core/n11067_2 ),
	.SUM(\top/processor/sha_core/n11067_1 )
);
defparam \top/processor/sha_core/n11067_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11066_s  (
	.I0(\top/processor/sha_core/h7 [22]),
	.I1(\top/processor/sha_core/h [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11067_2 ),
	.COUT(\top/processor/sha_core/n11066_2 ),
	.SUM(\top/processor/sha_core/n11066_1 )
);
defparam \top/processor/sha_core/n11066_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11065_s  (
	.I0(\top/processor/sha_core/h7 [23]),
	.I1(\top/processor/sha_core/h [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11066_2 ),
	.COUT(\top/processor/sha_core/n11065_2 ),
	.SUM(\top/processor/sha_core/n11065_1 )
);
defparam \top/processor/sha_core/n11065_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11064_s  (
	.I0(\top/processor/sha_core/h7 [24]),
	.I1(\top/processor/sha_core/h [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11065_2 ),
	.COUT(\top/processor/sha_core/n11064_2 ),
	.SUM(\top/processor/sha_core/n11064_1 )
);
defparam \top/processor/sha_core/n11064_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11063_s  (
	.I0(\top/processor/sha_core/h7 [25]),
	.I1(\top/processor/sha_core/h [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11064_2 ),
	.COUT(\top/processor/sha_core/n11063_2 ),
	.SUM(\top/processor/sha_core/n11063_1 )
);
defparam \top/processor/sha_core/n11063_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11062_s  (
	.I0(\top/processor/sha_core/h7 [26]),
	.I1(\top/processor/sha_core/h [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11063_2 ),
	.COUT(\top/processor/sha_core/n11062_2 ),
	.SUM(\top/processor/sha_core/n11062_1 )
);
defparam \top/processor/sha_core/n11062_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11061_s  (
	.I0(\top/processor/sha_core/h7 [27]),
	.I1(\top/processor/sha_core/h [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11062_2 ),
	.COUT(\top/processor/sha_core/n11061_2 ),
	.SUM(\top/processor/sha_core/n11061_1 )
);
defparam \top/processor/sha_core/n11061_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11060_s  (
	.I0(\top/processor/sha_core/h7 [28]),
	.I1(\top/processor/sha_core/h [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11061_2 ),
	.COUT(\top/processor/sha_core/n11060_2 ),
	.SUM(\top/processor/sha_core/n11060_1 )
);
defparam \top/processor/sha_core/n11060_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11059_s  (
	.I0(\top/processor/sha_core/h7 [29]),
	.I1(\top/processor/sha_core/h [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11060_2 ),
	.COUT(\top/processor/sha_core/n11059_2 ),
	.SUM(\top/processor/sha_core/n11059_1 )
);
defparam \top/processor/sha_core/n11059_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11058_s  (
	.I0(\top/processor/sha_core/h7 [30]),
	.I1(\top/processor/sha_core/h [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11059_2 ),
	.COUT(\top/processor/sha_core/n11058_2 ),
	.SUM(\top/processor/sha_core/n11058_1 )
);
defparam \top/processor/sha_core/n11058_s .ALU_MODE=0;
ALU \top/processor/sha_core/n11057_s  (
	.I0(\top/processor/sha_core/h7 [31]),
	.I1(\top/processor/sha_core/h [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n11058_2 ),
	.COUT(\top/processor/sha_core/n11057_0_COUT ),
	.SUM(\top/processor/sha_core/n11057_1 )
);
defparam \top/processor/sha_core/n11057_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10783_s  (
	.I0(\top/processor/sha_core/h [0]),
	.I1(\top/processor/sha_core/d [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10783_4 ),
	.SUM(\top/processor/sha_core/n10783_3 )
);
defparam \top/processor/sha_core/n10783_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10782_s  (
	.I0(\top/processor/sha_core/h [1]),
	.I1(\top/processor/sha_core/d [1]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10783_4 ),
	.COUT(\top/processor/sha_core/n10782_4 ),
	.SUM(\top/processor/sha_core/n10782_3 )
);
defparam \top/processor/sha_core/n10782_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10781_s  (
	.I0(\top/processor/sha_core/h [2]),
	.I1(\top/processor/sha_core/d [2]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10782_4 ),
	.COUT(\top/processor/sha_core/n10781_4 ),
	.SUM(\top/processor/sha_core/n10781_3 )
);
defparam \top/processor/sha_core/n10781_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10780_s  (
	.I0(\top/processor/sha_core/h [3]),
	.I1(\top/processor/sha_core/d [3]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10781_4 ),
	.COUT(\top/processor/sha_core/n10780_4 ),
	.SUM(\top/processor/sha_core/n10780_3 )
);
defparam \top/processor/sha_core/n10780_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10779_s  (
	.I0(\top/processor/sha_core/h [4]),
	.I1(\top/processor/sha_core/d [4]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10780_4 ),
	.COUT(\top/processor/sha_core/n10779_4 ),
	.SUM(\top/processor/sha_core/n10779_3 )
);
defparam \top/processor/sha_core/n10779_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10778_s  (
	.I0(\top/processor/sha_core/h [5]),
	.I1(\top/processor/sha_core/d [5]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10779_4 ),
	.COUT(\top/processor/sha_core/n10778_4 ),
	.SUM(\top/processor/sha_core/n10778_3 )
);
defparam \top/processor/sha_core/n10778_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10777_s  (
	.I0(\top/processor/sha_core/h [6]),
	.I1(\top/processor/sha_core/d [6]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10778_4 ),
	.COUT(\top/processor/sha_core/n10777_4 ),
	.SUM(\top/processor/sha_core/n10777_3 )
);
defparam \top/processor/sha_core/n10777_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10776_s  (
	.I0(\top/processor/sha_core/h [7]),
	.I1(\top/processor/sha_core/d [7]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10777_4 ),
	.COUT(\top/processor/sha_core/n10776_4 ),
	.SUM(\top/processor/sha_core/n10776_3 )
);
defparam \top/processor/sha_core/n10776_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10775_s  (
	.I0(\top/processor/sha_core/h [8]),
	.I1(\top/processor/sha_core/d [8]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10776_4 ),
	.COUT(\top/processor/sha_core/n10775_4 ),
	.SUM(\top/processor/sha_core/n10775_3 )
);
defparam \top/processor/sha_core/n10775_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10774_s  (
	.I0(\top/processor/sha_core/h [9]),
	.I1(\top/processor/sha_core/d [9]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10775_4 ),
	.COUT(\top/processor/sha_core/n10774_4 ),
	.SUM(\top/processor/sha_core/n10774_3 )
);
defparam \top/processor/sha_core/n10774_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10773_s  (
	.I0(\top/processor/sha_core/h [10]),
	.I1(\top/processor/sha_core/d [10]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10774_4 ),
	.COUT(\top/processor/sha_core/n10773_4 ),
	.SUM(\top/processor/sha_core/n10773_3 )
);
defparam \top/processor/sha_core/n10773_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10772_s  (
	.I0(\top/processor/sha_core/h [11]),
	.I1(\top/processor/sha_core/d [11]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10773_4 ),
	.COUT(\top/processor/sha_core/n10772_4 ),
	.SUM(\top/processor/sha_core/n10772_3 )
);
defparam \top/processor/sha_core/n10772_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10771_s  (
	.I0(\top/processor/sha_core/h [12]),
	.I1(\top/processor/sha_core/d [12]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10772_4 ),
	.COUT(\top/processor/sha_core/n10771_4 ),
	.SUM(\top/processor/sha_core/n10771_3 )
);
defparam \top/processor/sha_core/n10771_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10770_s  (
	.I0(\top/processor/sha_core/h [13]),
	.I1(\top/processor/sha_core/d [13]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10771_4 ),
	.COUT(\top/processor/sha_core/n10770_4 ),
	.SUM(\top/processor/sha_core/n10770_3 )
);
defparam \top/processor/sha_core/n10770_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10769_s  (
	.I0(\top/processor/sha_core/h [14]),
	.I1(\top/processor/sha_core/d [14]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10770_4 ),
	.COUT(\top/processor/sha_core/n10769_4 ),
	.SUM(\top/processor/sha_core/n10769_3 )
);
defparam \top/processor/sha_core/n10769_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10768_s  (
	.I0(\top/processor/sha_core/h [15]),
	.I1(\top/processor/sha_core/d [15]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10769_4 ),
	.COUT(\top/processor/sha_core/n10768_4 ),
	.SUM(\top/processor/sha_core/n10768_3 )
);
defparam \top/processor/sha_core/n10768_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10767_s  (
	.I0(\top/processor/sha_core/h [16]),
	.I1(\top/processor/sha_core/d [16]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10768_4 ),
	.COUT(\top/processor/sha_core/n10767_4 ),
	.SUM(\top/processor/sha_core/n10767_3 )
);
defparam \top/processor/sha_core/n10767_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10766_s  (
	.I0(\top/processor/sha_core/h [17]),
	.I1(\top/processor/sha_core/d [17]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10767_4 ),
	.COUT(\top/processor/sha_core/n10766_4 ),
	.SUM(\top/processor/sha_core/n10766_3 )
);
defparam \top/processor/sha_core/n10766_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10765_s  (
	.I0(\top/processor/sha_core/h [18]),
	.I1(\top/processor/sha_core/d [18]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10766_4 ),
	.COUT(\top/processor/sha_core/n10765_4 ),
	.SUM(\top/processor/sha_core/n10765_3 )
);
defparam \top/processor/sha_core/n10765_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10764_s  (
	.I0(\top/processor/sha_core/h [19]),
	.I1(\top/processor/sha_core/d [19]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10765_4 ),
	.COUT(\top/processor/sha_core/n10764_4 ),
	.SUM(\top/processor/sha_core/n10764_3 )
);
defparam \top/processor/sha_core/n10764_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10763_s  (
	.I0(\top/processor/sha_core/h [20]),
	.I1(\top/processor/sha_core/d [20]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10764_4 ),
	.COUT(\top/processor/sha_core/n10763_4 ),
	.SUM(\top/processor/sha_core/n10763_3 )
);
defparam \top/processor/sha_core/n10763_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10762_s  (
	.I0(\top/processor/sha_core/h [21]),
	.I1(\top/processor/sha_core/d [21]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10763_4 ),
	.COUT(\top/processor/sha_core/n10762_4 ),
	.SUM(\top/processor/sha_core/n10762_3 )
);
defparam \top/processor/sha_core/n10762_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10761_s  (
	.I0(\top/processor/sha_core/h [22]),
	.I1(\top/processor/sha_core/d [22]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10762_4 ),
	.COUT(\top/processor/sha_core/n10761_4 ),
	.SUM(\top/processor/sha_core/n10761_3 )
);
defparam \top/processor/sha_core/n10761_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10760_s  (
	.I0(\top/processor/sha_core/h [23]),
	.I1(\top/processor/sha_core/d [23]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10761_4 ),
	.COUT(\top/processor/sha_core/n10760_4 ),
	.SUM(\top/processor/sha_core/n10760_3 )
);
defparam \top/processor/sha_core/n10760_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10759_s  (
	.I0(\top/processor/sha_core/h [24]),
	.I1(\top/processor/sha_core/d [24]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10760_4 ),
	.COUT(\top/processor/sha_core/n10759_4 ),
	.SUM(\top/processor/sha_core/n10759_3 )
);
defparam \top/processor/sha_core/n10759_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10758_s  (
	.I0(\top/processor/sha_core/h [25]),
	.I1(\top/processor/sha_core/d [25]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10759_4 ),
	.COUT(\top/processor/sha_core/n10758_4 ),
	.SUM(\top/processor/sha_core/n10758_3 )
);
defparam \top/processor/sha_core/n10758_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10757_s  (
	.I0(\top/processor/sha_core/h [26]),
	.I1(\top/processor/sha_core/d [26]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10758_4 ),
	.COUT(\top/processor/sha_core/n10757_4 ),
	.SUM(\top/processor/sha_core/n10757_3 )
);
defparam \top/processor/sha_core/n10757_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10756_s  (
	.I0(\top/processor/sha_core/h [27]),
	.I1(\top/processor/sha_core/d [27]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10757_4 ),
	.COUT(\top/processor/sha_core/n10756_4 ),
	.SUM(\top/processor/sha_core/n10756_3 )
);
defparam \top/processor/sha_core/n10756_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10755_s  (
	.I0(\top/processor/sha_core/h [28]),
	.I1(\top/processor/sha_core/d [28]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10756_4 ),
	.COUT(\top/processor/sha_core/n10755_4 ),
	.SUM(\top/processor/sha_core/n10755_3 )
);
defparam \top/processor/sha_core/n10755_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10754_s  (
	.I0(\top/processor/sha_core/h [29]),
	.I1(\top/processor/sha_core/d [29]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10755_4 ),
	.COUT(\top/processor/sha_core/n10754_4 ),
	.SUM(\top/processor/sha_core/n10754_3 )
);
defparam \top/processor/sha_core/n10754_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10753_s  (
	.I0(\top/processor/sha_core/h [30]),
	.I1(\top/processor/sha_core/d [30]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10754_4 ),
	.COUT(\top/processor/sha_core/n10753_4 ),
	.SUM(\top/processor/sha_core/n10753_3 )
);
defparam \top/processor/sha_core/n10753_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10752_s  (
	.I0(\top/processor/sha_core/h [31]),
	.I1(\top/processor/sha_core/d [31]),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10753_4 ),
	.COUT(\top/processor/sha_core/n10752_0_COUT ),
	.SUM(\top/processor/sha_core/n10752_3 )
);
defparam \top/processor/sha_core/n10752_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10783_s0  (
	.I0(\top/processor/sha_core/n36_3 ),
	.I1(\top/processor/sha_core/n197_3 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10783_6 ),
	.SUM(\top/processor/sha_core/n10783_5 )
);
defparam \top/processor/sha_core/n10783_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10782_s0  (
	.I0(\top/processor/sha_core/n37_3 ),
	.I1(\top/processor/sha_core/n198_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10783_6 ),
	.COUT(\top/processor/sha_core/n10782_6 ),
	.SUM(\top/processor/sha_core/n10782_5 )
);
defparam \top/processor/sha_core/n10782_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10781_s0  (
	.I0(\top/processor/sha_core/n38_3 ),
	.I1(\top/processor/sha_core/n199_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10782_6 ),
	.COUT(\top/processor/sha_core/n10781_6 ),
	.SUM(\top/processor/sha_core/n10781_5 )
);
defparam \top/processor/sha_core/n10781_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10780_s0  (
	.I0(\top/processor/sha_core/n39_3 ),
	.I1(\top/processor/sha_core/n200_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10781_6 ),
	.COUT(\top/processor/sha_core/n10780_6 ),
	.SUM(\top/processor/sha_core/n10780_5 )
);
defparam \top/processor/sha_core/n10780_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10779_s0  (
	.I0(\top/processor/sha_core/n40_3 ),
	.I1(\top/processor/sha_core/n201_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10780_6 ),
	.COUT(\top/processor/sha_core/n10779_6 ),
	.SUM(\top/processor/sha_core/n10779_5 )
);
defparam \top/processor/sha_core/n10779_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10778_s0  (
	.I0(\top/processor/sha_core/n41_3 ),
	.I1(\top/processor/sha_core/n202_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10779_6 ),
	.COUT(\top/processor/sha_core/n10778_6 ),
	.SUM(\top/processor/sha_core/n10778_5 )
);
defparam \top/processor/sha_core/n10778_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10777_s0  (
	.I0(\top/processor/sha_core/n42_3 ),
	.I1(\top/processor/sha_core/n203_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10778_6 ),
	.COUT(\top/processor/sha_core/n10777_6 ),
	.SUM(\top/processor/sha_core/n10777_5 )
);
defparam \top/processor/sha_core/n10777_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10776_s0  (
	.I0(\top/processor/sha_core/n43_3 ),
	.I1(\top/processor/sha_core/n204_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10777_6 ),
	.COUT(\top/processor/sha_core/n10776_6 ),
	.SUM(\top/processor/sha_core/n10776_5 )
);
defparam \top/processor/sha_core/n10776_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10775_s0  (
	.I0(\top/processor/sha_core/n44_3 ),
	.I1(\top/processor/sha_core/n205_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10776_6 ),
	.COUT(\top/processor/sha_core/n10775_6 ),
	.SUM(\top/processor/sha_core/n10775_5 )
);
defparam \top/processor/sha_core/n10775_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10774_s0  (
	.I0(\top/processor/sha_core/n45_3 ),
	.I1(\top/processor/sha_core/n206_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10775_6 ),
	.COUT(\top/processor/sha_core/n10774_6 ),
	.SUM(\top/processor/sha_core/n10774_5 )
);
defparam \top/processor/sha_core/n10774_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10773_s0  (
	.I0(\top/processor/sha_core/n46_3 ),
	.I1(\top/processor/sha_core/n207_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10774_6 ),
	.COUT(\top/processor/sha_core/n10773_6 ),
	.SUM(\top/processor/sha_core/n10773_5 )
);
defparam \top/processor/sha_core/n10773_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10772_s0  (
	.I0(\top/processor/sha_core/n47_3 ),
	.I1(\top/processor/sha_core/n208_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10773_6 ),
	.COUT(\top/processor/sha_core/n10772_6 ),
	.SUM(\top/processor/sha_core/n10772_5 )
);
defparam \top/processor/sha_core/n10772_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10771_s0  (
	.I0(\top/processor/sha_core/n48_3 ),
	.I1(\top/processor/sha_core/n209_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10772_6 ),
	.COUT(\top/processor/sha_core/n10771_6 ),
	.SUM(\top/processor/sha_core/n10771_5 )
);
defparam \top/processor/sha_core/n10771_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10770_s0  (
	.I0(\top/processor/sha_core/n49_3 ),
	.I1(\top/processor/sha_core/n210_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10771_6 ),
	.COUT(\top/processor/sha_core/n10770_6 ),
	.SUM(\top/processor/sha_core/n10770_5 )
);
defparam \top/processor/sha_core/n10770_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10769_s0  (
	.I0(\top/processor/sha_core/n50_3 ),
	.I1(\top/processor/sha_core/n211_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10770_6 ),
	.COUT(\top/processor/sha_core/n10769_6 ),
	.SUM(\top/processor/sha_core/n10769_5 )
);
defparam \top/processor/sha_core/n10769_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10768_s0  (
	.I0(\top/processor/sha_core/n51_3 ),
	.I1(\top/processor/sha_core/n212_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10769_6 ),
	.COUT(\top/processor/sha_core/n10768_6 ),
	.SUM(\top/processor/sha_core/n10768_5 )
);
defparam \top/processor/sha_core/n10768_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10767_s0  (
	.I0(\top/processor/sha_core/n52_3 ),
	.I1(\top/processor/sha_core/n213_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10768_6 ),
	.COUT(\top/processor/sha_core/n10767_6 ),
	.SUM(\top/processor/sha_core/n10767_5 )
);
defparam \top/processor/sha_core/n10767_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10766_s0  (
	.I0(\top/processor/sha_core/n53_3 ),
	.I1(\top/processor/sha_core/n214_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10767_6 ),
	.COUT(\top/processor/sha_core/n10766_6 ),
	.SUM(\top/processor/sha_core/n10766_5 )
);
defparam \top/processor/sha_core/n10766_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10765_s0  (
	.I0(\top/processor/sha_core/n54_3 ),
	.I1(\top/processor/sha_core/n215_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10766_6 ),
	.COUT(\top/processor/sha_core/n10765_6 ),
	.SUM(\top/processor/sha_core/n10765_5 )
);
defparam \top/processor/sha_core/n10765_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10764_s0  (
	.I0(\top/processor/sha_core/n55_3 ),
	.I1(\top/processor/sha_core/n216_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10765_6 ),
	.COUT(\top/processor/sha_core/n10764_6 ),
	.SUM(\top/processor/sha_core/n10764_5 )
);
defparam \top/processor/sha_core/n10764_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10763_s0  (
	.I0(\top/processor/sha_core/n56_3 ),
	.I1(\top/processor/sha_core/n217_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10764_6 ),
	.COUT(\top/processor/sha_core/n10763_6 ),
	.SUM(\top/processor/sha_core/n10763_5 )
);
defparam \top/processor/sha_core/n10763_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10762_s0  (
	.I0(\top/processor/sha_core/n57_3 ),
	.I1(\top/processor/sha_core/n218_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10763_6 ),
	.COUT(\top/processor/sha_core/n10762_6 ),
	.SUM(\top/processor/sha_core/n10762_5 )
);
defparam \top/processor/sha_core/n10762_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10761_s0  (
	.I0(\top/processor/sha_core/n58_3 ),
	.I1(\top/processor/sha_core/n219_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10762_6 ),
	.COUT(\top/processor/sha_core/n10761_6 ),
	.SUM(\top/processor/sha_core/n10761_5 )
);
defparam \top/processor/sha_core/n10761_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10760_s0  (
	.I0(\top/processor/sha_core/n59_3 ),
	.I1(\top/processor/sha_core/n220_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10761_6 ),
	.COUT(\top/processor/sha_core/n10760_6 ),
	.SUM(\top/processor/sha_core/n10760_5 )
);
defparam \top/processor/sha_core/n10760_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10759_s0  (
	.I0(\top/processor/sha_core/n60_3 ),
	.I1(\top/processor/sha_core/n221_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10760_6 ),
	.COUT(\top/processor/sha_core/n10759_6 ),
	.SUM(\top/processor/sha_core/n10759_5 )
);
defparam \top/processor/sha_core/n10759_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10758_s0  (
	.I0(\top/processor/sha_core/n61_3 ),
	.I1(\top/processor/sha_core/n222_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10759_6 ),
	.COUT(\top/processor/sha_core/n10758_6 ),
	.SUM(\top/processor/sha_core/n10758_5 )
);
defparam \top/processor/sha_core/n10758_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10757_s0  (
	.I0(\top/processor/sha_core/n62_3 ),
	.I1(\top/processor/sha_core/n223_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10758_6 ),
	.COUT(\top/processor/sha_core/n10757_6 ),
	.SUM(\top/processor/sha_core/n10757_5 )
);
defparam \top/processor/sha_core/n10757_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10756_s0  (
	.I0(\top/processor/sha_core/n63_3 ),
	.I1(\top/processor/sha_core/n224_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10757_6 ),
	.COUT(\top/processor/sha_core/n10756_6 ),
	.SUM(\top/processor/sha_core/n10756_5 )
);
defparam \top/processor/sha_core/n10756_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10755_s0  (
	.I0(\top/processor/sha_core/n64_3 ),
	.I1(\top/processor/sha_core/n225_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10756_6 ),
	.COUT(\top/processor/sha_core/n10755_6 ),
	.SUM(\top/processor/sha_core/n10755_5 )
);
defparam \top/processor/sha_core/n10755_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10754_s0  (
	.I0(\top/processor/sha_core/n65_3 ),
	.I1(\top/processor/sha_core/n226_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10755_6 ),
	.COUT(\top/processor/sha_core/n10754_6 ),
	.SUM(\top/processor/sha_core/n10754_5 )
);
defparam \top/processor/sha_core/n10754_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10753_s0  (
	.I0(\top/processor/sha_core/n66_3 ),
	.I1(\top/processor/sha_core/n227_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10754_6 ),
	.COUT(\top/processor/sha_core/n10753_6 ),
	.SUM(\top/processor/sha_core/n10753_5 )
);
defparam \top/processor/sha_core/n10753_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10752_s0  (
	.I0(\top/processor/sha_core/n67_3 ),
	.I1(\top/processor/sha_core/n228_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10753_6 ),
	.COUT(\top/processor/sha_core/n10752_1_COUT ),
	.SUM(\top/processor/sha_core/n10752_5 )
);
defparam \top/processor/sha_core/n10752_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10783_s1  (
	.I0(\top/processor/sha_core/n293_7162 ),
	.I1(\top/processor/sha_core/n358_225 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10783_8 ),
	.SUM(\top/processor/sha_core/n10783_7 )
);
defparam \top/processor/sha_core/n10783_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10782_s1  (
	.I0(\top/processor/sha_core/n293_7164 ),
	.I1(\top/processor/sha_core/n357_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10783_8 ),
	.COUT(\top/processor/sha_core/n10782_8 ),
	.SUM(\top/processor/sha_core/n10782_7 )
);
defparam \top/processor/sha_core/n10782_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10781_s1  (
	.I0(\top/processor/sha_core/n293_7166 ),
	.I1(\top/processor/sha_core/n356_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10782_8 ),
	.COUT(\top/processor/sha_core/n10781_8 ),
	.SUM(\top/processor/sha_core/n10781_7 )
);
defparam \top/processor/sha_core/n10781_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10780_s1  (
	.I0(\top/processor/sha_core/n293_7168 ),
	.I1(\top/processor/sha_core/n355_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10781_8 ),
	.COUT(\top/processor/sha_core/n10780_8 ),
	.SUM(\top/processor/sha_core/n10780_7 )
);
defparam \top/processor/sha_core/n10780_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10779_s1  (
	.I0(\top/processor/sha_core/n293_7170 ),
	.I1(\top/processor/sha_core/n354_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10780_8 ),
	.COUT(\top/processor/sha_core/n10779_8 ),
	.SUM(\top/processor/sha_core/n10779_7 )
);
defparam \top/processor/sha_core/n10779_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10778_s1  (
	.I0(\top/processor/sha_core/n293_7172 ),
	.I1(\top/processor/sha_core/n353_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10779_8 ),
	.COUT(\top/processor/sha_core/n10778_8 ),
	.SUM(\top/processor/sha_core/n10778_7 )
);
defparam \top/processor/sha_core/n10778_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10777_s1  (
	.I0(\top/processor/sha_core/n293_7174 ),
	.I1(\top/processor/sha_core/n352_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10778_8 ),
	.COUT(\top/processor/sha_core/n10777_8 ),
	.SUM(\top/processor/sha_core/n10777_7 )
);
defparam \top/processor/sha_core/n10777_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10776_s1  (
	.I0(\top/processor/sha_core/n293_7176 ),
	.I1(\top/processor/sha_core/n351_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10777_8 ),
	.COUT(\top/processor/sha_core/n10776_8 ),
	.SUM(\top/processor/sha_core/n10776_7 )
);
defparam \top/processor/sha_core/n10776_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10775_s1  (
	.I0(\top/processor/sha_core/n293_7178 ),
	.I1(\top/processor/sha_core/n350_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10776_8 ),
	.COUT(\top/processor/sha_core/n10775_8 ),
	.SUM(\top/processor/sha_core/n10775_7 )
);
defparam \top/processor/sha_core/n10775_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10774_s1  (
	.I0(\top/processor/sha_core/n293_7180 ),
	.I1(\top/processor/sha_core/n349_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10775_8 ),
	.COUT(\top/processor/sha_core/n10774_8 ),
	.SUM(\top/processor/sha_core/n10774_7 )
);
defparam \top/processor/sha_core/n10774_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10773_s1  (
	.I0(\top/processor/sha_core/n293_7182 ),
	.I1(\top/processor/sha_core/n348_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10774_8 ),
	.COUT(\top/processor/sha_core/n10773_8 ),
	.SUM(\top/processor/sha_core/n10773_7 )
);
defparam \top/processor/sha_core/n10773_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10772_s1  (
	.I0(\top/processor/sha_core/n293_7184 ),
	.I1(\top/processor/sha_core/n347_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10773_8 ),
	.COUT(\top/processor/sha_core/n10772_8 ),
	.SUM(\top/processor/sha_core/n10772_7 )
);
defparam \top/processor/sha_core/n10772_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10771_s1  (
	.I0(\top/processor/sha_core/n293_7186 ),
	.I1(\top/processor/sha_core/n346_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10772_8 ),
	.COUT(\top/processor/sha_core/n10771_8 ),
	.SUM(\top/processor/sha_core/n10771_7 )
);
defparam \top/processor/sha_core/n10771_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10770_s1  (
	.I0(\top/processor/sha_core/n293_7188 ),
	.I1(\top/processor/sha_core/n345_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10771_8 ),
	.COUT(\top/processor/sha_core/n10770_8 ),
	.SUM(\top/processor/sha_core/n10770_7 )
);
defparam \top/processor/sha_core/n10770_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10769_s1  (
	.I0(\top/processor/sha_core/n293_7190 ),
	.I1(\top/processor/sha_core/n344_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10770_8 ),
	.COUT(\top/processor/sha_core/n10769_8 ),
	.SUM(\top/processor/sha_core/n10769_7 )
);
defparam \top/processor/sha_core/n10769_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10768_s1  (
	.I0(\top/processor/sha_core/n293_7192 ),
	.I1(\top/processor/sha_core/n343_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10769_8 ),
	.COUT(\top/processor/sha_core/n10768_8 ),
	.SUM(\top/processor/sha_core/n10768_7 )
);
defparam \top/processor/sha_core/n10768_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10767_s1  (
	.I0(\top/processor/sha_core/n293_7194 ),
	.I1(\top/processor/sha_core/n342_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10768_8 ),
	.COUT(\top/processor/sha_core/n10767_8 ),
	.SUM(\top/processor/sha_core/n10767_7 )
);
defparam \top/processor/sha_core/n10767_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10766_s1  (
	.I0(\top/processor/sha_core/n293_7196 ),
	.I1(\top/processor/sha_core/n341_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10767_8 ),
	.COUT(\top/processor/sha_core/n10766_8 ),
	.SUM(\top/processor/sha_core/n10766_7 )
);
defparam \top/processor/sha_core/n10766_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10765_s1  (
	.I0(\top/processor/sha_core/n293_7198 ),
	.I1(\top/processor/sha_core/n340_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10766_8 ),
	.COUT(\top/processor/sha_core/n10765_8 ),
	.SUM(\top/processor/sha_core/n10765_7 )
);
defparam \top/processor/sha_core/n10765_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10764_s1  (
	.I0(\top/processor/sha_core/n293_7200 ),
	.I1(\top/processor/sha_core/n339_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10765_8 ),
	.COUT(\top/processor/sha_core/n10764_8 ),
	.SUM(\top/processor/sha_core/n10764_7 )
);
defparam \top/processor/sha_core/n10764_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10763_s1  (
	.I0(\top/processor/sha_core/n293_7202 ),
	.I1(\top/processor/sha_core/n338_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10764_8 ),
	.COUT(\top/processor/sha_core/n10763_8 ),
	.SUM(\top/processor/sha_core/n10763_7 )
);
defparam \top/processor/sha_core/n10763_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10762_s1  (
	.I0(\top/processor/sha_core/n293_7204 ),
	.I1(\top/processor/sha_core/n337_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10763_8 ),
	.COUT(\top/processor/sha_core/n10762_8 ),
	.SUM(\top/processor/sha_core/n10762_7 )
);
defparam \top/processor/sha_core/n10762_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10761_s1  (
	.I0(\top/processor/sha_core/n293_7206 ),
	.I1(\top/processor/sha_core/n336_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10762_8 ),
	.COUT(\top/processor/sha_core/n10761_8 ),
	.SUM(\top/processor/sha_core/n10761_7 )
);
defparam \top/processor/sha_core/n10761_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10760_s1  (
	.I0(\top/processor/sha_core/n293_7208 ),
	.I1(\top/processor/sha_core/n335_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10761_8 ),
	.COUT(\top/processor/sha_core/n10760_8 ),
	.SUM(\top/processor/sha_core/n10760_7 )
);
defparam \top/processor/sha_core/n10760_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10759_s1  (
	.I0(\top/processor/sha_core/n293_7210 ),
	.I1(\top/processor/sha_core/n334_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10760_8 ),
	.COUT(\top/processor/sha_core/n10759_8 ),
	.SUM(\top/processor/sha_core/n10759_7 )
);
defparam \top/processor/sha_core/n10759_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10758_s1  (
	.I0(\top/processor/sha_core/n293_7212 ),
	.I1(\top/processor/sha_core/n333_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10759_8 ),
	.COUT(\top/processor/sha_core/n10758_8 ),
	.SUM(\top/processor/sha_core/n10758_7 )
);
defparam \top/processor/sha_core/n10758_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10757_s1  (
	.I0(\top/processor/sha_core/n293_7214 ),
	.I1(\top/processor/sha_core/n332_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10758_8 ),
	.COUT(\top/processor/sha_core/n10757_8 ),
	.SUM(\top/processor/sha_core/n10757_7 )
);
defparam \top/processor/sha_core/n10757_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10756_s1  (
	.I0(\top/processor/sha_core/n293_7216 ),
	.I1(\top/processor/sha_core/n331_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10757_8 ),
	.COUT(\top/processor/sha_core/n10756_8 ),
	.SUM(\top/processor/sha_core/n10756_7 )
);
defparam \top/processor/sha_core/n10756_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10755_s1  (
	.I0(\top/processor/sha_core/n293_7218 ),
	.I1(\top/processor/sha_core/n330_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10756_8 ),
	.COUT(\top/processor/sha_core/n10755_8 ),
	.SUM(\top/processor/sha_core/n10755_7 )
);
defparam \top/processor/sha_core/n10755_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10754_s1  (
	.I0(\top/processor/sha_core/n293_7220 ),
	.I1(\top/processor/sha_core/n329_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10755_8 ),
	.COUT(\top/processor/sha_core/n10754_8 ),
	.SUM(\top/processor/sha_core/n10754_7 )
);
defparam \top/processor/sha_core/n10754_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10753_s1  (
	.I0(\top/processor/sha_core/n293_7222 ),
	.I1(\top/processor/sha_core/n328_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10754_8 ),
	.COUT(\top/processor/sha_core/n10753_8 ),
	.SUM(\top/processor/sha_core/n10753_7 )
);
defparam \top/processor/sha_core/n10753_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10752_s1  (
	.I0(\top/processor/sha_core/n293_7224 ),
	.I1(\top/processor/sha_core/n327_225 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10753_8 ),
	.COUT(\top/processor/sha_core/n10752_2_COUT ),
	.SUM(\top/processor/sha_core/n10752_7 )
);
defparam \top/processor/sha_core/n10752_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10783_s2  (
	.I0(\top/processor/sha_core/n10783_3 ),
	.I1(\top/processor/sha_core/n10783_5 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10783_10 ),
	.SUM(\top/processor/sha_core/n10783_9 )
);
defparam \top/processor/sha_core/n10783_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10782_s2  (
	.I0(\top/processor/sha_core/n10782_3 ),
	.I1(\top/processor/sha_core/n10782_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10783_10 ),
	.COUT(\top/processor/sha_core/n10782_10 ),
	.SUM(\top/processor/sha_core/n10782_9 )
);
defparam \top/processor/sha_core/n10782_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10781_s2  (
	.I0(\top/processor/sha_core/n10781_3 ),
	.I1(\top/processor/sha_core/n10781_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10782_10 ),
	.COUT(\top/processor/sha_core/n10781_10 ),
	.SUM(\top/processor/sha_core/n10781_9 )
);
defparam \top/processor/sha_core/n10781_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10780_s2  (
	.I0(\top/processor/sha_core/n10780_3 ),
	.I1(\top/processor/sha_core/n10780_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10781_10 ),
	.COUT(\top/processor/sha_core/n10780_10 ),
	.SUM(\top/processor/sha_core/n10780_9 )
);
defparam \top/processor/sha_core/n10780_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10779_s2  (
	.I0(\top/processor/sha_core/n10779_3 ),
	.I1(\top/processor/sha_core/n10779_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10780_10 ),
	.COUT(\top/processor/sha_core/n10779_10 ),
	.SUM(\top/processor/sha_core/n10779_9 )
);
defparam \top/processor/sha_core/n10779_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10778_s2  (
	.I0(\top/processor/sha_core/n10778_3 ),
	.I1(\top/processor/sha_core/n10778_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10779_10 ),
	.COUT(\top/processor/sha_core/n10778_10 ),
	.SUM(\top/processor/sha_core/n10778_9 )
);
defparam \top/processor/sha_core/n10778_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10777_s2  (
	.I0(\top/processor/sha_core/n10777_3 ),
	.I1(\top/processor/sha_core/n10777_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10778_10 ),
	.COUT(\top/processor/sha_core/n10777_10 ),
	.SUM(\top/processor/sha_core/n10777_9 )
);
defparam \top/processor/sha_core/n10777_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10776_s2  (
	.I0(\top/processor/sha_core/n10776_3 ),
	.I1(\top/processor/sha_core/n10776_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10777_10 ),
	.COUT(\top/processor/sha_core/n10776_10 ),
	.SUM(\top/processor/sha_core/n10776_9 )
);
defparam \top/processor/sha_core/n10776_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10775_s2  (
	.I0(\top/processor/sha_core/n10775_3 ),
	.I1(\top/processor/sha_core/n10775_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10776_10 ),
	.COUT(\top/processor/sha_core/n10775_10 ),
	.SUM(\top/processor/sha_core/n10775_9 )
);
defparam \top/processor/sha_core/n10775_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10774_s2  (
	.I0(\top/processor/sha_core/n10774_3 ),
	.I1(\top/processor/sha_core/n10774_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10775_10 ),
	.COUT(\top/processor/sha_core/n10774_10 ),
	.SUM(\top/processor/sha_core/n10774_9 )
);
defparam \top/processor/sha_core/n10774_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10773_s2  (
	.I0(\top/processor/sha_core/n10773_3 ),
	.I1(\top/processor/sha_core/n10773_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10774_10 ),
	.COUT(\top/processor/sha_core/n10773_10 ),
	.SUM(\top/processor/sha_core/n10773_9 )
);
defparam \top/processor/sha_core/n10773_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10772_s2  (
	.I0(\top/processor/sha_core/n10772_3 ),
	.I1(\top/processor/sha_core/n10772_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10773_10 ),
	.COUT(\top/processor/sha_core/n10772_10 ),
	.SUM(\top/processor/sha_core/n10772_9 )
);
defparam \top/processor/sha_core/n10772_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10771_s2  (
	.I0(\top/processor/sha_core/n10771_3 ),
	.I1(\top/processor/sha_core/n10771_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10772_10 ),
	.COUT(\top/processor/sha_core/n10771_10 ),
	.SUM(\top/processor/sha_core/n10771_9 )
);
defparam \top/processor/sha_core/n10771_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10770_s2  (
	.I0(\top/processor/sha_core/n10770_3 ),
	.I1(\top/processor/sha_core/n10770_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10771_10 ),
	.COUT(\top/processor/sha_core/n10770_10 ),
	.SUM(\top/processor/sha_core/n10770_9 )
);
defparam \top/processor/sha_core/n10770_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10769_s2  (
	.I0(\top/processor/sha_core/n10769_3 ),
	.I1(\top/processor/sha_core/n10769_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10770_10 ),
	.COUT(\top/processor/sha_core/n10769_10 ),
	.SUM(\top/processor/sha_core/n10769_9 )
);
defparam \top/processor/sha_core/n10769_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10768_s2  (
	.I0(\top/processor/sha_core/n10768_3 ),
	.I1(\top/processor/sha_core/n10768_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10769_10 ),
	.COUT(\top/processor/sha_core/n10768_10 ),
	.SUM(\top/processor/sha_core/n10768_9 )
);
defparam \top/processor/sha_core/n10768_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10767_s2  (
	.I0(\top/processor/sha_core/n10767_3 ),
	.I1(\top/processor/sha_core/n10767_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10768_10 ),
	.COUT(\top/processor/sha_core/n10767_10 ),
	.SUM(\top/processor/sha_core/n10767_9 )
);
defparam \top/processor/sha_core/n10767_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10766_s2  (
	.I0(\top/processor/sha_core/n10766_3 ),
	.I1(\top/processor/sha_core/n10766_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10767_10 ),
	.COUT(\top/processor/sha_core/n10766_10 ),
	.SUM(\top/processor/sha_core/n10766_9 )
);
defparam \top/processor/sha_core/n10766_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10765_s2  (
	.I0(\top/processor/sha_core/n10765_3 ),
	.I1(\top/processor/sha_core/n10765_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10766_10 ),
	.COUT(\top/processor/sha_core/n10765_10 ),
	.SUM(\top/processor/sha_core/n10765_9 )
);
defparam \top/processor/sha_core/n10765_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10764_s2  (
	.I0(\top/processor/sha_core/n10764_3 ),
	.I1(\top/processor/sha_core/n10764_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10765_10 ),
	.COUT(\top/processor/sha_core/n10764_10 ),
	.SUM(\top/processor/sha_core/n10764_9 )
);
defparam \top/processor/sha_core/n10764_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10763_s2  (
	.I0(\top/processor/sha_core/n10763_3 ),
	.I1(\top/processor/sha_core/n10763_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10764_10 ),
	.COUT(\top/processor/sha_core/n10763_10 ),
	.SUM(\top/processor/sha_core/n10763_9 )
);
defparam \top/processor/sha_core/n10763_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10762_s2  (
	.I0(\top/processor/sha_core/n10762_3 ),
	.I1(\top/processor/sha_core/n10762_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10763_10 ),
	.COUT(\top/processor/sha_core/n10762_10 ),
	.SUM(\top/processor/sha_core/n10762_9 )
);
defparam \top/processor/sha_core/n10762_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10761_s2  (
	.I0(\top/processor/sha_core/n10761_3 ),
	.I1(\top/processor/sha_core/n10761_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10762_10 ),
	.COUT(\top/processor/sha_core/n10761_10 ),
	.SUM(\top/processor/sha_core/n10761_9 )
);
defparam \top/processor/sha_core/n10761_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10760_s2  (
	.I0(\top/processor/sha_core/n10760_3 ),
	.I1(\top/processor/sha_core/n10760_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10761_10 ),
	.COUT(\top/processor/sha_core/n10760_10 ),
	.SUM(\top/processor/sha_core/n10760_9 )
);
defparam \top/processor/sha_core/n10760_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10759_s2  (
	.I0(\top/processor/sha_core/n10759_3 ),
	.I1(\top/processor/sha_core/n10759_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10760_10 ),
	.COUT(\top/processor/sha_core/n10759_10 ),
	.SUM(\top/processor/sha_core/n10759_9 )
);
defparam \top/processor/sha_core/n10759_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10758_s2  (
	.I0(\top/processor/sha_core/n10758_3 ),
	.I1(\top/processor/sha_core/n10758_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10759_10 ),
	.COUT(\top/processor/sha_core/n10758_10 ),
	.SUM(\top/processor/sha_core/n10758_9 )
);
defparam \top/processor/sha_core/n10758_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10757_s2  (
	.I0(\top/processor/sha_core/n10757_3 ),
	.I1(\top/processor/sha_core/n10757_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10758_10 ),
	.COUT(\top/processor/sha_core/n10757_10 ),
	.SUM(\top/processor/sha_core/n10757_9 )
);
defparam \top/processor/sha_core/n10757_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10756_s2  (
	.I0(\top/processor/sha_core/n10756_3 ),
	.I1(\top/processor/sha_core/n10756_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10757_10 ),
	.COUT(\top/processor/sha_core/n10756_10 ),
	.SUM(\top/processor/sha_core/n10756_9 )
);
defparam \top/processor/sha_core/n10756_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10755_s2  (
	.I0(\top/processor/sha_core/n10755_3 ),
	.I1(\top/processor/sha_core/n10755_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10756_10 ),
	.COUT(\top/processor/sha_core/n10755_10 ),
	.SUM(\top/processor/sha_core/n10755_9 )
);
defparam \top/processor/sha_core/n10755_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10754_s2  (
	.I0(\top/processor/sha_core/n10754_3 ),
	.I1(\top/processor/sha_core/n10754_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10755_10 ),
	.COUT(\top/processor/sha_core/n10754_10 ),
	.SUM(\top/processor/sha_core/n10754_9 )
);
defparam \top/processor/sha_core/n10754_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10753_s2  (
	.I0(\top/processor/sha_core/n10753_3 ),
	.I1(\top/processor/sha_core/n10753_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10754_10 ),
	.COUT(\top/processor/sha_core/n10753_10 ),
	.SUM(\top/processor/sha_core/n10753_9 )
);
defparam \top/processor/sha_core/n10753_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10752_s2  (
	.I0(\top/processor/sha_core/n10752_3 ),
	.I1(\top/processor/sha_core/n10752_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10753_10 ),
	.COUT(\top/processor/sha_core/n10752_3_COUT ),
	.SUM(\top/processor/sha_core/n10752_9 )
);
defparam \top/processor/sha_core/n10752_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10783_s3  (
	.I0(\top/processor/sha_core/n10783_9 ),
	.I1(\top/processor/sha_core/n10783_7 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10783_12 ),
	.SUM(\top/processor/sha_core/n10783_11 )
);
defparam \top/processor/sha_core/n10783_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10782_s3  (
	.I0(\top/processor/sha_core/n10782_9 ),
	.I1(\top/processor/sha_core/n10782_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10783_12 ),
	.COUT(\top/processor/sha_core/n10782_12 ),
	.SUM(\top/processor/sha_core/n10782_11 )
);
defparam \top/processor/sha_core/n10782_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10781_s3  (
	.I0(\top/processor/sha_core/n10781_9 ),
	.I1(\top/processor/sha_core/n10781_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10782_12 ),
	.COUT(\top/processor/sha_core/n10781_12 ),
	.SUM(\top/processor/sha_core/n10781_11 )
);
defparam \top/processor/sha_core/n10781_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10780_s3  (
	.I0(\top/processor/sha_core/n10780_9 ),
	.I1(\top/processor/sha_core/n10780_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10781_12 ),
	.COUT(\top/processor/sha_core/n10780_12 ),
	.SUM(\top/processor/sha_core/n10780_11 )
);
defparam \top/processor/sha_core/n10780_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10779_s3  (
	.I0(\top/processor/sha_core/n10779_9 ),
	.I1(\top/processor/sha_core/n10779_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10780_12 ),
	.COUT(\top/processor/sha_core/n10779_12 ),
	.SUM(\top/processor/sha_core/n10779_11 )
);
defparam \top/processor/sha_core/n10779_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10778_s3  (
	.I0(\top/processor/sha_core/n10778_9 ),
	.I1(\top/processor/sha_core/n10778_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10779_12 ),
	.COUT(\top/processor/sha_core/n10778_12 ),
	.SUM(\top/processor/sha_core/n10778_11 )
);
defparam \top/processor/sha_core/n10778_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10777_s3  (
	.I0(\top/processor/sha_core/n10777_9 ),
	.I1(\top/processor/sha_core/n10777_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10778_12 ),
	.COUT(\top/processor/sha_core/n10777_12 ),
	.SUM(\top/processor/sha_core/n10777_11 )
);
defparam \top/processor/sha_core/n10777_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10776_s3  (
	.I0(\top/processor/sha_core/n10776_9 ),
	.I1(\top/processor/sha_core/n10776_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10777_12 ),
	.COUT(\top/processor/sha_core/n10776_12 ),
	.SUM(\top/processor/sha_core/n10776_11 )
);
defparam \top/processor/sha_core/n10776_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10775_s3  (
	.I0(\top/processor/sha_core/n10775_9 ),
	.I1(\top/processor/sha_core/n10775_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10776_12 ),
	.COUT(\top/processor/sha_core/n10775_12 ),
	.SUM(\top/processor/sha_core/n10775_11 )
);
defparam \top/processor/sha_core/n10775_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10774_s3  (
	.I0(\top/processor/sha_core/n10774_9 ),
	.I1(\top/processor/sha_core/n10774_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10775_12 ),
	.COUT(\top/processor/sha_core/n10774_12 ),
	.SUM(\top/processor/sha_core/n10774_11 )
);
defparam \top/processor/sha_core/n10774_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10773_s3  (
	.I0(\top/processor/sha_core/n10773_9 ),
	.I1(\top/processor/sha_core/n10773_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10774_12 ),
	.COUT(\top/processor/sha_core/n10773_12 ),
	.SUM(\top/processor/sha_core/n10773_11 )
);
defparam \top/processor/sha_core/n10773_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10772_s3  (
	.I0(\top/processor/sha_core/n10772_9 ),
	.I1(\top/processor/sha_core/n10772_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10773_12 ),
	.COUT(\top/processor/sha_core/n10772_12 ),
	.SUM(\top/processor/sha_core/n10772_11 )
);
defparam \top/processor/sha_core/n10772_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10771_s3  (
	.I0(\top/processor/sha_core/n10771_9 ),
	.I1(\top/processor/sha_core/n10771_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10772_12 ),
	.COUT(\top/processor/sha_core/n10771_12 ),
	.SUM(\top/processor/sha_core/n10771_11 )
);
defparam \top/processor/sha_core/n10771_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10770_s3  (
	.I0(\top/processor/sha_core/n10770_9 ),
	.I1(\top/processor/sha_core/n10770_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10771_12 ),
	.COUT(\top/processor/sha_core/n10770_12 ),
	.SUM(\top/processor/sha_core/n10770_11 )
);
defparam \top/processor/sha_core/n10770_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10769_s3  (
	.I0(\top/processor/sha_core/n10769_9 ),
	.I1(\top/processor/sha_core/n10769_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10770_12 ),
	.COUT(\top/processor/sha_core/n10769_12 ),
	.SUM(\top/processor/sha_core/n10769_11 )
);
defparam \top/processor/sha_core/n10769_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10768_s3  (
	.I0(\top/processor/sha_core/n10768_9 ),
	.I1(\top/processor/sha_core/n10768_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10769_12 ),
	.COUT(\top/processor/sha_core/n10768_12 ),
	.SUM(\top/processor/sha_core/n10768_11 )
);
defparam \top/processor/sha_core/n10768_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10767_s3  (
	.I0(\top/processor/sha_core/n10767_9 ),
	.I1(\top/processor/sha_core/n10767_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10768_12 ),
	.COUT(\top/processor/sha_core/n10767_12 ),
	.SUM(\top/processor/sha_core/n10767_11 )
);
defparam \top/processor/sha_core/n10767_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10766_s3  (
	.I0(\top/processor/sha_core/n10766_9 ),
	.I1(\top/processor/sha_core/n10766_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10767_12 ),
	.COUT(\top/processor/sha_core/n10766_12 ),
	.SUM(\top/processor/sha_core/n10766_11 )
);
defparam \top/processor/sha_core/n10766_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10765_s3  (
	.I0(\top/processor/sha_core/n10765_9 ),
	.I1(\top/processor/sha_core/n10765_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10766_12 ),
	.COUT(\top/processor/sha_core/n10765_12 ),
	.SUM(\top/processor/sha_core/n10765_11 )
);
defparam \top/processor/sha_core/n10765_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10764_s3  (
	.I0(\top/processor/sha_core/n10764_9 ),
	.I1(\top/processor/sha_core/n10764_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10765_12 ),
	.COUT(\top/processor/sha_core/n10764_12 ),
	.SUM(\top/processor/sha_core/n10764_11 )
);
defparam \top/processor/sha_core/n10764_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10763_s3  (
	.I0(\top/processor/sha_core/n10763_9 ),
	.I1(\top/processor/sha_core/n10763_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10764_12 ),
	.COUT(\top/processor/sha_core/n10763_12 ),
	.SUM(\top/processor/sha_core/n10763_11 )
);
defparam \top/processor/sha_core/n10763_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10762_s3  (
	.I0(\top/processor/sha_core/n10762_9 ),
	.I1(\top/processor/sha_core/n10762_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10763_12 ),
	.COUT(\top/processor/sha_core/n10762_12 ),
	.SUM(\top/processor/sha_core/n10762_11 )
);
defparam \top/processor/sha_core/n10762_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10761_s3  (
	.I0(\top/processor/sha_core/n10761_9 ),
	.I1(\top/processor/sha_core/n10761_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10762_12 ),
	.COUT(\top/processor/sha_core/n10761_12 ),
	.SUM(\top/processor/sha_core/n10761_11 )
);
defparam \top/processor/sha_core/n10761_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10760_s3  (
	.I0(\top/processor/sha_core/n10760_9 ),
	.I1(\top/processor/sha_core/n10760_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10761_12 ),
	.COUT(\top/processor/sha_core/n10760_12 ),
	.SUM(\top/processor/sha_core/n10760_11 )
);
defparam \top/processor/sha_core/n10760_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10759_s3  (
	.I0(\top/processor/sha_core/n10759_9 ),
	.I1(\top/processor/sha_core/n10759_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10760_12 ),
	.COUT(\top/processor/sha_core/n10759_12 ),
	.SUM(\top/processor/sha_core/n10759_11 )
);
defparam \top/processor/sha_core/n10759_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10758_s3  (
	.I0(\top/processor/sha_core/n10758_9 ),
	.I1(\top/processor/sha_core/n10758_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10759_12 ),
	.COUT(\top/processor/sha_core/n10758_12 ),
	.SUM(\top/processor/sha_core/n10758_11 )
);
defparam \top/processor/sha_core/n10758_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10757_s3  (
	.I0(\top/processor/sha_core/n10757_9 ),
	.I1(\top/processor/sha_core/n10757_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10758_12 ),
	.COUT(\top/processor/sha_core/n10757_12 ),
	.SUM(\top/processor/sha_core/n10757_11 )
);
defparam \top/processor/sha_core/n10757_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10756_s3  (
	.I0(\top/processor/sha_core/n10756_9 ),
	.I1(\top/processor/sha_core/n10756_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10757_12 ),
	.COUT(\top/processor/sha_core/n10756_12 ),
	.SUM(\top/processor/sha_core/n10756_11 )
);
defparam \top/processor/sha_core/n10756_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10755_s3  (
	.I0(\top/processor/sha_core/n10755_9 ),
	.I1(\top/processor/sha_core/n10755_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10756_12 ),
	.COUT(\top/processor/sha_core/n10755_12 ),
	.SUM(\top/processor/sha_core/n10755_11 )
);
defparam \top/processor/sha_core/n10755_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10754_s3  (
	.I0(\top/processor/sha_core/n10754_9 ),
	.I1(\top/processor/sha_core/n10754_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10755_12 ),
	.COUT(\top/processor/sha_core/n10754_12 ),
	.SUM(\top/processor/sha_core/n10754_11 )
);
defparam \top/processor/sha_core/n10754_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10753_s3  (
	.I0(\top/processor/sha_core/n10753_9 ),
	.I1(\top/processor/sha_core/n10753_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10754_12 ),
	.COUT(\top/processor/sha_core/n10753_12 ),
	.SUM(\top/processor/sha_core/n10753_11 )
);
defparam \top/processor/sha_core/n10753_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10752_s3  (
	.I0(\top/processor/sha_core/n10752_9 ),
	.I1(\top/processor/sha_core/n10752_7 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10753_12 ),
	.COUT(\top/processor/sha_core/n10752_4_COUT ),
	.SUM(\top/processor/sha_core/n10752_11 )
);
defparam \top/processor/sha_core/n10752_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10816_s  (
	.I0(\top/processor/sha_core/h [0]),
	.I1(\top/processor/sha_core/n36_3 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10816_4 ),
	.SUM(\top/processor/sha_core/n10816_3 )
);
defparam \top/processor/sha_core/n10816_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10815_s  (
	.I0(\top/processor/sha_core/h [1]),
	.I1(\top/processor/sha_core/n37_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10816_4 ),
	.COUT(\top/processor/sha_core/n10815_4 ),
	.SUM(\top/processor/sha_core/n10815_3 )
);
defparam \top/processor/sha_core/n10815_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10814_s  (
	.I0(\top/processor/sha_core/h [2]),
	.I1(\top/processor/sha_core/n38_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10815_4 ),
	.COUT(\top/processor/sha_core/n10814_4 ),
	.SUM(\top/processor/sha_core/n10814_3 )
);
defparam \top/processor/sha_core/n10814_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10813_s  (
	.I0(\top/processor/sha_core/h [3]),
	.I1(\top/processor/sha_core/n39_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10814_4 ),
	.COUT(\top/processor/sha_core/n10813_4 ),
	.SUM(\top/processor/sha_core/n10813_3 )
);
defparam \top/processor/sha_core/n10813_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10812_s  (
	.I0(\top/processor/sha_core/h [4]),
	.I1(\top/processor/sha_core/n40_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10813_4 ),
	.COUT(\top/processor/sha_core/n10812_4 ),
	.SUM(\top/processor/sha_core/n10812_3 )
);
defparam \top/processor/sha_core/n10812_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10811_s  (
	.I0(\top/processor/sha_core/h [5]),
	.I1(\top/processor/sha_core/n41_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10812_4 ),
	.COUT(\top/processor/sha_core/n10811_4 ),
	.SUM(\top/processor/sha_core/n10811_3 )
);
defparam \top/processor/sha_core/n10811_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10810_s  (
	.I0(\top/processor/sha_core/h [6]),
	.I1(\top/processor/sha_core/n42_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10811_4 ),
	.COUT(\top/processor/sha_core/n10810_4 ),
	.SUM(\top/processor/sha_core/n10810_3 )
);
defparam \top/processor/sha_core/n10810_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10809_s  (
	.I0(\top/processor/sha_core/h [7]),
	.I1(\top/processor/sha_core/n43_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10810_4 ),
	.COUT(\top/processor/sha_core/n10809_4 ),
	.SUM(\top/processor/sha_core/n10809_3 )
);
defparam \top/processor/sha_core/n10809_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10808_s  (
	.I0(\top/processor/sha_core/h [8]),
	.I1(\top/processor/sha_core/n44_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10809_4 ),
	.COUT(\top/processor/sha_core/n10808_4 ),
	.SUM(\top/processor/sha_core/n10808_3 )
);
defparam \top/processor/sha_core/n10808_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10807_s  (
	.I0(\top/processor/sha_core/h [9]),
	.I1(\top/processor/sha_core/n45_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10808_4 ),
	.COUT(\top/processor/sha_core/n10807_4 ),
	.SUM(\top/processor/sha_core/n10807_3 )
);
defparam \top/processor/sha_core/n10807_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10806_s  (
	.I0(\top/processor/sha_core/h [10]),
	.I1(\top/processor/sha_core/n46_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10807_4 ),
	.COUT(\top/processor/sha_core/n10806_4 ),
	.SUM(\top/processor/sha_core/n10806_3 )
);
defparam \top/processor/sha_core/n10806_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10805_s  (
	.I0(\top/processor/sha_core/h [11]),
	.I1(\top/processor/sha_core/n47_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10806_4 ),
	.COUT(\top/processor/sha_core/n10805_4 ),
	.SUM(\top/processor/sha_core/n10805_3 )
);
defparam \top/processor/sha_core/n10805_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10804_s  (
	.I0(\top/processor/sha_core/h [12]),
	.I1(\top/processor/sha_core/n48_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10805_4 ),
	.COUT(\top/processor/sha_core/n10804_4 ),
	.SUM(\top/processor/sha_core/n10804_3 )
);
defparam \top/processor/sha_core/n10804_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10803_s  (
	.I0(\top/processor/sha_core/h [13]),
	.I1(\top/processor/sha_core/n49_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10804_4 ),
	.COUT(\top/processor/sha_core/n10803_4 ),
	.SUM(\top/processor/sha_core/n10803_3 )
);
defparam \top/processor/sha_core/n10803_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10802_s  (
	.I0(\top/processor/sha_core/h [14]),
	.I1(\top/processor/sha_core/n50_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10803_4 ),
	.COUT(\top/processor/sha_core/n10802_4 ),
	.SUM(\top/processor/sha_core/n10802_3 )
);
defparam \top/processor/sha_core/n10802_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10801_s  (
	.I0(\top/processor/sha_core/h [15]),
	.I1(\top/processor/sha_core/n51_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10802_4 ),
	.COUT(\top/processor/sha_core/n10801_4 ),
	.SUM(\top/processor/sha_core/n10801_3 )
);
defparam \top/processor/sha_core/n10801_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10800_s  (
	.I0(\top/processor/sha_core/h [16]),
	.I1(\top/processor/sha_core/n52_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10801_4 ),
	.COUT(\top/processor/sha_core/n10800_4 ),
	.SUM(\top/processor/sha_core/n10800_3 )
);
defparam \top/processor/sha_core/n10800_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10799_s  (
	.I0(\top/processor/sha_core/h [17]),
	.I1(\top/processor/sha_core/n53_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10800_4 ),
	.COUT(\top/processor/sha_core/n10799_4 ),
	.SUM(\top/processor/sha_core/n10799_3 )
);
defparam \top/processor/sha_core/n10799_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10798_s  (
	.I0(\top/processor/sha_core/h [18]),
	.I1(\top/processor/sha_core/n54_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10799_4 ),
	.COUT(\top/processor/sha_core/n10798_4 ),
	.SUM(\top/processor/sha_core/n10798_3 )
);
defparam \top/processor/sha_core/n10798_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10797_s  (
	.I0(\top/processor/sha_core/h [19]),
	.I1(\top/processor/sha_core/n55_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10798_4 ),
	.COUT(\top/processor/sha_core/n10797_4 ),
	.SUM(\top/processor/sha_core/n10797_3 )
);
defparam \top/processor/sha_core/n10797_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10796_s  (
	.I0(\top/processor/sha_core/h [20]),
	.I1(\top/processor/sha_core/n56_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10797_4 ),
	.COUT(\top/processor/sha_core/n10796_4 ),
	.SUM(\top/processor/sha_core/n10796_3 )
);
defparam \top/processor/sha_core/n10796_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10795_s  (
	.I0(\top/processor/sha_core/h [21]),
	.I1(\top/processor/sha_core/n57_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10796_4 ),
	.COUT(\top/processor/sha_core/n10795_4 ),
	.SUM(\top/processor/sha_core/n10795_3 )
);
defparam \top/processor/sha_core/n10795_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10794_s  (
	.I0(\top/processor/sha_core/h [22]),
	.I1(\top/processor/sha_core/n58_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10795_4 ),
	.COUT(\top/processor/sha_core/n10794_4 ),
	.SUM(\top/processor/sha_core/n10794_3 )
);
defparam \top/processor/sha_core/n10794_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10793_s  (
	.I0(\top/processor/sha_core/h [23]),
	.I1(\top/processor/sha_core/n59_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10794_4 ),
	.COUT(\top/processor/sha_core/n10793_4 ),
	.SUM(\top/processor/sha_core/n10793_3 )
);
defparam \top/processor/sha_core/n10793_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10792_s  (
	.I0(\top/processor/sha_core/h [24]),
	.I1(\top/processor/sha_core/n60_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10793_4 ),
	.COUT(\top/processor/sha_core/n10792_4 ),
	.SUM(\top/processor/sha_core/n10792_3 )
);
defparam \top/processor/sha_core/n10792_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10791_s  (
	.I0(\top/processor/sha_core/h [25]),
	.I1(\top/processor/sha_core/n61_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10792_4 ),
	.COUT(\top/processor/sha_core/n10791_4 ),
	.SUM(\top/processor/sha_core/n10791_3 )
);
defparam \top/processor/sha_core/n10791_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10790_s  (
	.I0(\top/processor/sha_core/h [26]),
	.I1(\top/processor/sha_core/n62_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10791_4 ),
	.COUT(\top/processor/sha_core/n10790_4 ),
	.SUM(\top/processor/sha_core/n10790_3 )
);
defparam \top/processor/sha_core/n10790_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10789_s  (
	.I0(\top/processor/sha_core/h [27]),
	.I1(\top/processor/sha_core/n63_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10790_4 ),
	.COUT(\top/processor/sha_core/n10789_4 ),
	.SUM(\top/processor/sha_core/n10789_3 )
);
defparam \top/processor/sha_core/n10789_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10788_s  (
	.I0(\top/processor/sha_core/h [28]),
	.I1(\top/processor/sha_core/n64_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10789_4 ),
	.COUT(\top/processor/sha_core/n10788_4 ),
	.SUM(\top/processor/sha_core/n10788_3 )
);
defparam \top/processor/sha_core/n10788_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10787_s  (
	.I0(\top/processor/sha_core/h [29]),
	.I1(\top/processor/sha_core/n65_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10788_4 ),
	.COUT(\top/processor/sha_core/n10787_4 ),
	.SUM(\top/processor/sha_core/n10787_3 )
);
defparam \top/processor/sha_core/n10787_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10786_s  (
	.I0(\top/processor/sha_core/h [30]),
	.I1(\top/processor/sha_core/n66_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10787_4 ),
	.COUT(\top/processor/sha_core/n10786_4 ),
	.SUM(\top/processor/sha_core/n10786_3 )
);
defparam \top/processor/sha_core/n10786_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10785_s  (
	.I0(\top/processor/sha_core/h [31]),
	.I1(\top/processor/sha_core/n67_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10786_4 ),
	.COUT(\top/processor/sha_core/n10785_0_COUT ),
	.SUM(\top/processor/sha_core/n10785_3 )
);
defparam \top/processor/sha_core/n10785_s .ALU_MODE=0;
ALU \top/processor/sha_core/n10816_s0  (
	.I0(\top/processor/sha_core/n197_3 ),
	.I1(\top/processor/sha_core/n293_7162 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10816_6 ),
	.SUM(\top/processor/sha_core/n10816_5 )
);
defparam \top/processor/sha_core/n10816_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10815_s0  (
	.I0(\top/processor/sha_core/n198_3 ),
	.I1(\top/processor/sha_core/n293_7164 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10816_6 ),
	.COUT(\top/processor/sha_core/n10815_6 ),
	.SUM(\top/processor/sha_core/n10815_5 )
);
defparam \top/processor/sha_core/n10815_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10814_s0  (
	.I0(\top/processor/sha_core/n199_3 ),
	.I1(\top/processor/sha_core/n293_7166 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10815_6 ),
	.COUT(\top/processor/sha_core/n10814_6 ),
	.SUM(\top/processor/sha_core/n10814_5 )
);
defparam \top/processor/sha_core/n10814_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10813_s0  (
	.I0(\top/processor/sha_core/n200_3 ),
	.I1(\top/processor/sha_core/n293_7168 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10814_6 ),
	.COUT(\top/processor/sha_core/n10813_6 ),
	.SUM(\top/processor/sha_core/n10813_5 )
);
defparam \top/processor/sha_core/n10813_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10812_s0  (
	.I0(\top/processor/sha_core/n201_3 ),
	.I1(\top/processor/sha_core/n293_7170 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10813_6 ),
	.COUT(\top/processor/sha_core/n10812_6 ),
	.SUM(\top/processor/sha_core/n10812_5 )
);
defparam \top/processor/sha_core/n10812_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10811_s0  (
	.I0(\top/processor/sha_core/n202_3 ),
	.I1(\top/processor/sha_core/n293_7172 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10812_6 ),
	.COUT(\top/processor/sha_core/n10811_6 ),
	.SUM(\top/processor/sha_core/n10811_5 )
);
defparam \top/processor/sha_core/n10811_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10810_s0  (
	.I0(\top/processor/sha_core/n203_3 ),
	.I1(\top/processor/sha_core/n293_7174 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10811_6 ),
	.COUT(\top/processor/sha_core/n10810_6 ),
	.SUM(\top/processor/sha_core/n10810_5 )
);
defparam \top/processor/sha_core/n10810_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10809_s0  (
	.I0(\top/processor/sha_core/n204_3 ),
	.I1(\top/processor/sha_core/n293_7176 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10810_6 ),
	.COUT(\top/processor/sha_core/n10809_6 ),
	.SUM(\top/processor/sha_core/n10809_5 )
);
defparam \top/processor/sha_core/n10809_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10808_s0  (
	.I0(\top/processor/sha_core/n205_3 ),
	.I1(\top/processor/sha_core/n293_7178 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10809_6 ),
	.COUT(\top/processor/sha_core/n10808_6 ),
	.SUM(\top/processor/sha_core/n10808_5 )
);
defparam \top/processor/sha_core/n10808_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10807_s0  (
	.I0(\top/processor/sha_core/n206_3 ),
	.I1(\top/processor/sha_core/n293_7180 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10808_6 ),
	.COUT(\top/processor/sha_core/n10807_6 ),
	.SUM(\top/processor/sha_core/n10807_5 )
);
defparam \top/processor/sha_core/n10807_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10806_s0  (
	.I0(\top/processor/sha_core/n207_3 ),
	.I1(\top/processor/sha_core/n293_7182 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10807_6 ),
	.COUT(\top/processor/sha_core/n10806_6 ),
	.SUM(\top/processor/sha_core/n10806_5 )
);
defparam \top/processor/sha_core/n10806_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10805_s0  (
	.I0(\top/processor/sha_core/n208_3 ),
	.I1(\top/processor/sha_core/n293_7184 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10806_6 ),
	.COUT(\top/processor/sha_core/n10805_6 ),
	.SUM(\top/processor/sha_core/n10805_5 )
);
defparam \top/processor/sha_core/n10805_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10804_s0  (
	.I0(\top/processor/sha_core/n209_3 ),
	.I1(\top/processor/sha_core/n293_7186 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10805_6 ),
	.COUT(\top/processor/sha_core/n10804_6 ),
	.SUM(\top/processor/sha_core/n10804_5 )
);
defparam \top/processor/sha_core/n10804_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10803_s0  (
	.I0(\top/processor/sha_core/n210_3 ),
	.I1(\top/processor/sha_core/n293_7188 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10804_6 ),
	.COUT(\top/processor/sha_core/n10803_6 ),
	.SUM(\top/processor/sha_core/n10803_5 )
);
defparam \top/processor/sha_core/n10803_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10802_s0  (
	.I0(\top/processor/sha_core/n211_3 ),
	.I1(\top/processor/sha_core/n293_7190 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10803_6 ),
	.COUT(\top/processor/sha_core/n10802_6 ),
	.SUM(\top/processor/sha_core/n10802_5 )
);
defparam \top/processor/sha_core/n10802_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10801_s0  (
	.I0(\top/processor/sha_core/n212_3 ),
	.I1(\top/processor/sha_core/n293_7192 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10802_6 ),
	.COUT(\top/processor/sha_core/n10801_6 ),
	.SUM(\top/processor/sha_core/n10801_5 )
);
defparam \top/processor/sha_core/n10801_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10800_s0  (
	.I0(\top/processor/sha_core/n213_3 ),
	.I1(\top/processor/sha_core/n293_7194 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10801_6 ),
	.COUT(\top/processor/sha_core/n10800_6 ),
	.SUM(\top/processor/sha_core/n10800_5 )
);
defparam \top/processor/sha_core/n10800_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10799_s0  (
	.I0(\top/processor/sha_core/n214_3 ),
	.I1(\top/processor/sha_core/n293_7196 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10800_6 ),
	.COUT(\top/processor/sha_core/n10799_6 ),
	.SUM(\top/processor/sha_core/n10799_5 )
);
defparam \top/processor/sha_core/n10799_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10798_s0  (
	.I0(\top/processor/sha_core/n215_3 ),
	.I1(\top/processor/sha_core/n293_7198 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10799_6 ),
	.COUT(\top/processor/sha_core/n10798_6 ),
	.SUM(\top/processor/sha_core/n10798_5 )
);
defparam \top/processor/sha_core/n10798_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10797_s0  (
	.I0(\top/processor/sha_core/n216_3 ),
	.I1(\top/processor/sha_core/n293_7200 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10798_6 ),
	.COUT(\top/processor/sha_core/n10797_6 ),
	.SUM(\top/processor/sha_core/n10797_5 )
);
defparam \top/processor/sha_core/n10797_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10796_s0  (
	.I0(\top/processor/sha_core/n217_3 ),
	.I1(\top/processor/sha_core/n293_7202 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10797_6 ),
	.COUT(\top/processor/sha_core/n10796_6 ),
	.SUM(\top/processor/sha_core/n10796_5 )
);
defparam \top/processor/sha_core/n10796_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10795_s0  (
	.I0(\top/processor/sha_core/n218_3 ),
	.I1(\top/processor/sha_core/n293_7204 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10796_6 ),
	.COUT(\top/processor/sha_core/n10795_6 ),
	.SUM(\top/processor/sha_core/n10795_5 )
);
defparam \top/processor/sha_core/n10795_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10794_s0  (
	.I0(\top/processor/sha_core/n219_3 ),
	.I1(\top/processor/sha_core/n293_7206 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10795_6 ),
	.COUT(\top/processor/sha_core/n10794_6 ),
	.SUM(\top/processor/sha_core/n10794_5 )
);
defparam \top/processor/sha_core/n10794_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10793_s0  (
	.I0(\top/processor/sha_core/n220_3 ),
	.I1(\top/processor/sha_core/n293_7208 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10794_6 ),
	.COUT(\top/processor/sha_core/n10793_6 ),
	.SUM(\top/processor/sha_core/n10793_5 )
);
defparam \top/processor/sha_core/n10793_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10792_s0  (
	.I0(\top/processor/sha_core/n221_3 ),
	.I1(\top/processor/sha_core/n293_7210 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10793_6 ),
	.COUT(\top/processor/sha_core/n10792_6 ),
	.SUM(\top/processor/sha_core/n10792_5 )
);
defparam \top/processor/sha_core/n10792_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10791_s0  (
	.I0(\top/processor/sha_core/n222_3 ),
	.I1(\top/processor/sha_core/n293_7212 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10792_6 ),
	.COUT(\top/processor/sha_core/n10791_6 ),
	.SUM(\top/processor/sha_core/n10791_5 )
);
defparam \top/processor/sha_core/n10791_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10790_s0  (
	.I0(\top/processor/sha_core/n223_3 ),
	.I1(\top/processor/sha_core/n293_7214 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10791_6 ),
	.COUT(\top/processor/sha_core/n10790_6 ),
	.SUM(\top/processor/sha_core/n10790_5 )
);
defparam \top/processor/sha_core/n10790_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10789_s0  (
	.I0(\top/processor/sha_core/n224_3 ),
	.I1(\top/processor/sha_core/n293_7216 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10790_6 ),
	.COUT(\top/processor/sha_core/n10789_6 ),
	.SUM(\top/processor/sha_core/n10789_5 )
);
defparam \top/processor/sha_core/n10789_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10788_s0  (
	.I0(\top/processor/sha_core/n225_3 ),
	.I1(\top/processor/sha_core/n293_7218 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10789_6 ),
	.COUT(\top/processor/sha_core/n10788_6 ),
	.SUM(\top/processor/sha_core/n10788_5 )
);
defparam \top/processor/sha_core/n10788_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10787_s0  (
	.I0(\top/processor/sha_core/n226_3 ),
	.I1(\top/processor/sha_core/n293_7220 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10788_6 ),
	.COUT(\top/processor/sha_core/n10787_6 ),
	.SUM(\top/processor/sha_core/n10787_5 )
);
defparam \top/processor/sha_core/n10787_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10786_s0  (
	.I0(\top/processor/sha_core/n227_3 ),
	.I1(\top/processor/sha_core/n293_7222 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10787_6 ),
	.COUT(\top/processor/sha_core/n10786_6 ),
	.SUM(\top/processor/sha_core/n10786_5 )
);
defparam \top/processor/sha_core/n10786_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10785_s0  (
	.I0(\top/processor/sha_core/n228_3 ),
	.I1(\top/processor/sha_core/n293_7224 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10786_6 ),
	.COUT(\top/processor/sha_core/n10785_1_COUT ),
	.SUM(\top/processor/sha_core/n10785_5 )
);
defparam \top/processor/sha_core/n10785_s0 .ALU_MODE=0;
ALU \top/processor/sha_core/n10816_s1  (
	.I0(\top/processor/sha_core/n358_225 ),
	.I1(\top/processor/sha_core/n424_3 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10816_8 ),
	.SUM(\top/processor/sha_core/n10816_7 )
);
defparam \top/processor/sha_core/n10816_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10815_s1  (
	.I0(\top/processor/sha_core/n357_225 ),
	.I1(\top/processor/sha_core/n425_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10816_8 ),
	.COUT(\top/processor/sha_core/n10815_8 ),
	.SUM(\top/processor/sha_core/n10815_7 )
);
defparam \top/processor/sha_core/n10815_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10814_s1  (
	.I0(\top/processor/sha_core/n356_225 ),
	.I1(\top/processor/sha_core/n426_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10815_8 ),
	.COUT(\top/processor/sha_core/n10814_8 ),
	.SUM(\top/processor/sha_core/n10814_7 )
);
defparam \top/processor/sha_core/n10814_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10813_s1  (
	.I0(\top/processor/sha_core/n355_225 ),
	.I1(\top/processor/sha_core/n427_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10814_8 ),
	.COUT(\top/processor/sha_core/n10813_8 ),
	.SUM(\top/processor/sha_core/n10813_7 )
);
defparam \top/processor/sha_core/n10813_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10812_s1  (
	.I0(\top/processor/sha_core/n354_225 ),
	.I1(\top/processor/sha_core/n428_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10813_8 ),
	.COUT(\top/processor/sha_core/n10812_8 ),
	.SUM(\top/processor/sha_core/n10812_7 )
);
defparam \top/processor/sha_core/n10812_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10811_s1  (
	.I0(\top/processor/sha_core/n353_225 ),
	.I1(\top/processor/sha_core/n429_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10812_8 ),
	.COUT(\top/processor/sha_core/n10811_8 ),
	.SUM(\top/processor/sha_core/n10811_7 )
);
defparam \top/processor/sha_core/n10811_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10810_s1  (
	.I0(\top/processor/sha_core/n352_225 ),
	.I1(\top/processor/sha_core/n430_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10811_8 ),
	.COUT(\top/processor/sha_core/n10810_8 ),
	.SUM(\top/processor/sha_core/n10810_7 )
);
defparam \top/processor/sha_core/n10810_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10809_s1  (
	.I0(\top/processor/sha_core/n351_225 ),
	.I1(\top/processor/sha_core/n431_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10810_8 ),
	.COUT(\top/processor/sha_core/n10809_8 ),
	.SUM(\top/processor/sha_core/n10809_7 )
);
defparam \top/processor/sha_core/n10809_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10808_s1  (
	.I0(\top/processor/sha_core/n350_225 ),
	.I1(\top/processor/sha_core/n432_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10809_8 ),
	.COUT(\top/processor/sha_core/n10808_8 ),
	.SUM(\top/processor/sha_core/n10808_7 )
);
defparam \top/processor/sha_core/n10808_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10807_s1  (
	.I0(\top/processor/sha_core/n349_225 ),
	.I1(\top/processor/sha_core/n433_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10808_8 ),
	.COUT(\top/processor/sha_core/n10807_8 ),
	.SUM(\top/processor/sha_core/n10807_7 )
);
defparam \top/processor/sha_core/n10807_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10806_s1  (
	.I0(\top/processor/sha_core/n348_225 ),
	.I1(\top/processor/sha_core/n434_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10807_8 ),
	.COUT(\top/processor/sha_core/n10806_8 ),
	.SUM(\top/processor/sha_core/n10806_7 )
);
defparam \top/processor/sha_core/n10806_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10805_s1  (
	.I0(\top/processor/sha_core/n347_225 ),
	.I1(\top/processor/sha_core/n435_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10806_8 ),
	.COUT(\top/processor/sha_core/n10805_8 ),
	.SUM(\top/processor/sha_core/n10805_7 )
);
defparam \top/processor/sha_core/n10805_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10804_s1  (
	.I0(\top/processor/sha_core/n346_225 ),
	.I1(\top/processor/sha_core/n436_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10805_8 ),
	.COUT(\top/processor/sha_core/n10804_8 ),
	.SUM(\top/processor/sha_core/n10804_7 )
);
defparam \top/processor/sha_core/n10804_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10803_s1  (
	.I0(\top/processor/sha_core/n345_225 ),
	.I1(\top/processor/sha_core/n437_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10804_8 ),
	.COUT(\top/processor/sha_core/n10803_8 ),
	.SUM(\top/processor/sha_core/n10803_7 )
);
defparam \top/processor/sha_core/n10803_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10802_s1  (
	.I0(\top/processor/sha_core/n344_225 ),
	.I1(\top/processor/sha_core/n438_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10803_8 ),
	.COUT(\top/processor/sha_core/n10802_8 ),
	.SUM(\top/processor/sha_core/n10802_7 )
);
defparam \top/processor/sha_core/n10802_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10801_s1  (
	.I0(\top/processor/sha_core/n343_225 ),
	.I1(\top/processor/sha_core/n439_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10802_8 ),
	.COUT(\top/processor/sha_core/n10801_8 ),
	.SUM(\top/processor/sha_core/n10801_7 )
);
defparam \top/processor/sha_core/n10801_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10800_s1  (
	.I0(\top/processor/sha_core/n342_225 ),
	.I1(\top/processor/sha_core/n440_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10801_8 ),
	.COUT(\top/processor/sha_core/n10800_8 ),
	.SUM(\top/processor/sha_core/n10800_7 )
);
defparam \top/processor/sha_core/n10800_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10799_s1  (
	.I0(\top/processor/sha_core/n341_225 ),
	.I1(\top/processor/sha_core/n441_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10800_8 ),
	.COUT(\top/processor/sha_core/n10799_8 ),
	.SUM(\top/processor/sha_core/n10799_7 )
);
defparam \top/processor/sha_core/n10799_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10798_s1  (
	.I0(\top/processor/sha_core/n340_225 ),
	.I1(\top/processor/sha_core/n442_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10799_8 ),
	.COUT(\top/processor/sha_core/n10798_8 ),
	.SUM(\top/processor/sha_core/n10798_7 )
);
defparam \top/processor/sha_core/n10798_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10797_s1  (
	.I0(\top/processor/sha_core/n339_225 ),
	.I1(\top/processor/sha_core/n443_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10798_8 ),
	.COUT(\top/processor/sha_core/n10797_8 ),
	.SUM(\top/processor/sha_core/n10797_7 )
);
defparam \top/processor/sha_core/n10797_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10796_s1  (
	.I0(\top/processor/sha_core/n338_225 ),
	.I1(\top/processor/sha_core/n444_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10797_8 ),
	.COUT(\top/processor/sha_core/n10796_8 ),
	.SUM(\top/processor/sha_core/n10796_7 )
);
defparam \top/processor/sha_core/n10796_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10795_s1  (
	.I0(\top/processor/sha_core/n337_225 ),
	.I1(\top/processor/sha_core/n445_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10796_8 ),
	.COUT(\top/processor/sha_core/n10795_8 ),
	.SUM(\top/processor/sha_core/n10795_7 )
);
defparam \top/processor/sha_core/n10795_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10794_s1  (
	.I0(\top/processor/sha_core/n336_225 ),
	.I1(\top/processor/sha_core/n446_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10795_8 ),
	.COUT(\top/processor/sha_core/n10794_8 ),
	.SUM(\top/processor/sha_core/n10794_7 )
);
defparam \top/processor/sha_core/n10794_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10793_s1  (
	.I0(\top/processor/sha_core/n335_225 ),
	.I1(\top/processor/sha_core/n447_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10794_8 ),
	.COUT(\top/processor/sha_core/n10793_8 ),
	.SUM(\top/processor/sha_core/n10793_7 )
);
defparam \top/processor/sha_core/n10793_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10792_s1  (
	.I0(\top/processor/sha_core/n334_225 ),
	.I1(\top/processor/sha_core/n448_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10793_8 ),
	.COUT(\top/processor/sha_core/n10792_8 ),
	.SUM(\top/processor/sha_core/n10792_7 )
);
defparam \top/processor/sha_core/n10792_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10791_s1  (
	.I0(\top/processor/sha_core/n333_225 ),
	.I1(\top/processor/sha_core/n449_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10792_8 ),
	.COUT(\top/processor/sha_core/n10791_8 ),
	.SUM(\top/processor/sha_core/n10791_7 )
);
defparam \top/processor/sha_core/n10791_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10790_s1  (
	.I0(\top/processor/sha_core/n332_225 ),
	.I1(\top/processor/sha_core/n450_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10791_8 ),
	.COUT(\top/processor/sha_core/n10790_8 ),
	.SUM(\top/processor/sha_core/n10790_7 )
);
defparam \top/processor/sha_core/n10790_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10789_s1  (
	.I0(\top/processor/sha_core/n331_225 ),
	.I1(\top/processor/sha_core/n451_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10790_8 ),
	.COUT(\top/processor/sha_core/n10789_8 ),
	.SUM(\top/processor/sha_core/n10789_7 )
);
defparam \top/processor/sha_core/n10789_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10788_s1  (
	.I0(\top/processor/sha_core/n330_225 ),
	.I1(\top/processor/sha_core/n452_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10789_8 ),
	.COUT(\top/processor/sha_core/n10788_8 ),
	.SUM(\top/processor/sha_core/n10788_7 )
);
defparam \top/processor/sha_core/n10788_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10787_s1  (
	.I0(\top/processor/sha_core/n329_225 ),
	.I1(\top/processor/sha_core/n453_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10788_8 ),
	.COUT(\top/processor/sha_core/n10787_8 ),
	.SUM(\top/processor/sha_core/n10787_7 )
);
defparam \top/processor/sha_core/n10787_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10786_s1  (
	.I0(\top/processor/sha_core/n328_225 ),
	.I1(\top/processor/sha_core/n454_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10787_8 ),
	.COUT(\top/processor/sha_core/n10786_8 ),
	.SUM(\top/processor/sha_core/n10786_7 )
);
defparam \top/processor/sha_core/n10786_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10785_s1  (
	.I0(\top/processor/sha_core/n327_225 ),
	.I1(\top/processor/sha_core/n455_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10786_8 ),
	.COUT(\top/processor/sha_core/n10785_2_COUT ),
	.SUM(\top/processor/sha_core/n10785_7 )
);
defparam \top/processor/sha_core/n10785_s1 .ALU_MODE=0;
ALU \top/processor/sha_core/n10816_s2  (
	.I0(\top/processor/sha_core/n10816_3 ),
	.I1(\top/processor/sha_core/n10816_5 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10816_10 ),
	.SUM(\top/processor/sha_core/n10816_9 )
);
defparam \top/processor/sha_core/n10816_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10815_s2  (
	.I0(\top/processor/sha_core/n10815_3 ),
	.I1(\top/processor/sha_core/n10815_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10816_10 ),
	.COUT(\top/processor/sha_core/n10815_10 ),
	.SUM(\top/processor/sha_core/n10815_9 )
);
defparam \top/processor/sha_core/n10815_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10814_s2  (
	.I0(\top/processor/sha_core/n10814_3 ),
	.I1(\top/processor/sha_core/n10814_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10815_10 ),
	.COUT(\top/processor/sha_core/n10814_10 ),
	.SUM(\top/processor/sha_core/n10814_9 )
);
defparam \top/processor/sha_core/n10814_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10813_s2  (
	.I0(\top/processor/sha_core/n10813_3 ),
	.I1(\top/processor/sha_core/n10813_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10814_10 ),
	.COUT(\top/processor/sha_core/n10813_10 ),
	.SUM(\top/processor/sha_core/n10813_9 )
);
defparam \top/processor/sha_core/n10813_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10812_s2  (
	.I0(\top/processor/sha_core/n10812_3 ),
	.I1(\top/processor/sha_core/n10812_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10813_10 ),
	.COUT(\top/processor/sha_core/n10812_10 ),
	.SUM(\top/processor/sha_core/n10812_9 )
);
defparam \top/processor/sha_core/n10812_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10811_s2  (
	.I0(\top/processor/sha_core/n10811_3 ),
	.I1(\top/processor/sha_core/n10811_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10812_10 ),
	.COUT(\top/processor/sha_core/n10811_10 ),
	.SUM(\top/processor/sha_core/n10811_9 )
);
defparam \top/processor/sha_core/n10811_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10810_s2  (
	.I0(\top/processor/sha_core/n10810_3 ),
	.I1(\top/processor/sha_core/n10810_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10811_10 ),
	.COUT(\top/processor/sha_core/n10810_10 ),
	.SUM(\top/processor/sha_core/n10810_9 )
);
defparam \top/processor/sha_core/n10810_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10809_s2  (
	.I0(\top/processor/sha_core/n10809_3 ),
	.I1(\top/processor/sha_core/n10809_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10810_10 ),
	.COUT(\top/processor/sha_core/n10809_10 ),
	.SUM(\top/processor/sha_core/n10809_9 )
);
defparam \top/processor/sha_core/n10809_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10808_s2  (
	.I0(\top/processor/sha_core/n10808_3 ),
	.I1(\top/processor/sha_core/n10808_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10809_10 ),
	.COUT(\top/processor/sha_core/n10808_10 ),
	.SUM(\top/processor/sha_core/n10808_9 )
);
defparam \top/processor/sha_core/n10808_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10807_s2  (
	.I0(\top/processor/sha_core/n10807_3 ),
	.I1(\top/processor/sha_core/n10807_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10808_10 ),
	.COUT(\top/processor/sha_core/n10807_10 ),
	.SUM(\top/processor/sha_core/n10807_9 )
);
defparam \top/processor/sha_core/n10807_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10806_s2  (
	.I0(\top/processor/sha_core/n10806_3 ),
	.I1(\top/processor/sha_core/n10806_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10807_10 ),
	.COUT(\top/processor/sha_core/n10806_10 ),
	.SUM(\top/processor/sha_core/n10806_9 )
);
defparam \top/processor/sha_core/n10806_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10805_s2  (
	.I0(\top/processor/sha_core/n10805_3 ),
	.I1(\top/processor/sha_core/n10805_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10806_10 ),
	.COUT(\top/processor/sha_core/n10805_10 ),
	.SUM(\top/processor/sha_core/n10805_9 )
);
defparam \top/processor/sha_core/n10805_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10804_s2  (
	.I0(\top/processor/sha_core/n10804_3 ),
	.I1(\top/processor/sha_core/n10804_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10805_10 ),
	.COUT(\top/processor/sha_core/n10804_10 ),
	.SUM(\top/processor/sha_core/n10804_9 )
);
defparam \top/processor/sha_core/n10804_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10803_s2  (
	.I0(\top/processor/sha_core/n10803_3 ),
	.I1(\top/processor/sha_core/n10803_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10804_10 ),
	.COUT(\top/processor/sha_core/n10803_10 ),
	.SUM(\top/processor/sha_core/n10803_9 )
);
defparam \top/processor/sha_core/n10803_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10802_s2  (
	.I0(\top/processor/sha_core/n10802_3 ),
	.I1(\top/processor/sha_core/n10802_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10803_10 ),
	.COUT(\top/processor/sha_core/n10802_10 ),
	.SUM(\top/processor/sha_core/n10802_9 )
);
defparam \top/processor/sha_core/n10802_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10801_s2  (
	.I0(\top/processor/sha_core/n10801_3 ),
	.I1(\top/processor/sha_core/n10801_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10802_10 ),
	.COUT(\top/processor/sha_core/n10801_10 ),
	.SUM(\top/processor/sha_core/n10801_9 )
);
defparam \top/processor/sha_core/n10801_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10800_s2  (
	.I0(\top/processor/sha_core/n10800_3 ),
	.I1(\top/processor/sha_core/n10800_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10801_10 ),
	.COUT(\top/processor/sha_core/n10800_10 ),
	.SUM(\top/processor/sha_core/n10800_9 )
);
defparam \top/processor/sha_core/n10800_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10799_s2  (
	.I0(\top/processor/sha_core/n10799_3 ),
	.I1(\top/processor/sha_core/n10799_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10800_10 ),
	.COUT(\top/processor/sha_core/n10799_10 ),
	.SUM(\top/processor/sha_core/n10799_9 )
);
defparam \top/processor/sha_core/n10799_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10798_s2  (
	.I0(\top/processor/sha_core/n10798_3 ),
	.I1(\top/processor/sha_core/n10798_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10799_10 ),
	.COUT(\top/processor/sha_core/n10798_10 ),
	.SUM(\top/processor/sha_core/n10798_9 )
);
defparam \top/processor/sha_core/n10798_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10797_s2  (
	.I0(\top/processor/sha_core/n10797_3 ),
	.I1(\top/processor/sha_core/n10797_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10798_10 ),
	.COUT(\top/processor/sha_core/n10797_10 ),
	.SUM(\top/processor/sha_core/n10797_9 )
);
defparam \top/processor/sha_core/n10797_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10796_s2  (
	.I0(\top/processor/sha_core/n10796_3 ),
	.I1(\top/processor/sha_core/n10796_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10797_10 ),
	.COUT(\top/processor/sha_core/n10796_10 ),
	.SUM(\top/processor/sha_core/n10796_9 )
);
defparam \top/processor/sha_core/n10796_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10795_s2  (
	.I0(\top/processor/sha_core/n10795_3 ),
	.I1(\top/processor/sha_core/n10795_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10796_10 ),
	.COUT(\top/processor/sha_core/n10795_10 ),
	.SUM(\top/processor/sha_core/n10795_9 )
);
defparam \top/processor/sha_core/n10795_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10794_s2  (
	.I0(\top/processor/sha_core/n10794_3 ),
	.I1(\top/processor/sha_core/n10794_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10795_10 ),
	.COUT(\top/processor/sha_core/n10794_10 ),
	.SUM(\top/processor/sha_core/n10794_9 )
);
defparam \top/processor/sha_core/n10794_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10793_s2  (
	.I0(\top/processor/sha_core/n10793_3 ),
	.I1(\top/processor/sha_core/n10793_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10794_10 ),
	.COUT(\top/processor/sha_core/n10793_10 ),
	.SUM(\top/processor/sha_core/n10793_9 )
);
defparam \top/processor/sha_core/n10793_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10792_s2  (
	.I0(\top/processor/sha_core/n10792_3 ),
	.I1(\top/processor/sha_core/n10792_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10793_10 ),
	.COUT(\top/processor/sha_core/n10792_10 ),
	.SUM(\top/processor/sha_core/n10792_9 )
);
defparam \top/processor/sha_core/n10792_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10791_s2  (
	.I0(\top/processor/sha_core/n10791_3 ),
	.I1(\top/processor/sha_core/n10791_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10792_10 ),
	.COUT(\top/processor/sha_core/n10791_10 ),
	.SUM(\top/processor/sha_core/n10791_9 )
);
defparam \top/processor/sha_core/n10791_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10790_s2  (
	.I0(\top/processor/sha_core/n10790_3 ),
	.I1(\top/processor/sha_core/n10790_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10791_10 ),
	.COUT(\top/processor/sha_core/n10790_10 ),
	.SUM(\top/processor/sha_core/n10790_9 )
);
defparam \top/processor/sha_core/n10790_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10789_s2  (
	.I0(\top/processor/sha_core/n10789_3 ),
	.I1(\top/processor/sha_core/n10789_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10790_10 ),
	.COUT(\top/processor/sha_core/n10789_10 ),
	.SUM(\top/processor/sha_core/n10789_9 )
);
defparam \top/processor/sha_core/n10789_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10788_s2  (
	.I0(\top/processor/sha_core/n10788_3 ),
	.I1(\top/processor/sha_core/n10788_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10789_10 ),
	.COUT(\top/processor/sha_core/n10788_10 ),
	.SUM(\top/processor/sha_core/n10788_9 )
);
defparam \top/processor/sha_core/n10788_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10787_s2  (
	.I0(\top/processor/sha_core/n10787_3 ),
	.I1(\top/processor/sha_core/n10787_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10788_10 ),
	.COUT(\top/processor/sha_core/n10787_10 ),
	.SUM(\top/processor/sha_core/n10787_9 )
);
defparam \top/processor/sha_core/n10787_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10786_s2  (
	.I0(\top/processor/sha_core/n10786_3 ),
	.I1(\top/processor/sha_core/n10786_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10787_10 ),
	.COUT(\top/processor/sha_core/n10786_10 ),
	.SUM(\top/processor/sha_core/n10786_9 )
);
defparam \top/processor/sha_core/n10786_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10785_s2  (
	.I0(\top/processor/sha_core/n10785_3 ),
	.I1(\top/processor/sha_core/n10785_5 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10786_10 ),
	.COUT(\top/processor/sha_core/n10785_3_COUT ),
	.SUM(\top/processor/sha_core/n10785_9 )
);
defparam \top/processor/sha_core/n10785_s2 .ALU_MODE=0;
ALU \top/processor/sha_core/n10816_s3  (
	.I0(\top/processor/sha_core/n10816_7 ),
	.I1(\top/processor/sha_core/n584_3 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10816_12 ),
	.SUM(\top/processor/sha_core/n10816_11 )
);
defparam \top/processor/sha_core/n10816_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10815_s3  (
	.I0(\top/processor/sha_core/n10815_7 ),
	.I1(\top/processor/sha_core/n585_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10816_12 ),
	.COUT(\top/processor/sha_core/n10815_12 ),
	.SUM(\top/processor/sha_core/n10815_11 )
);
defparam \top/processor/sha_core/n10815_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10814_s3  (
	.I0(\top/processor/sha_core/n10814_7 ),
	.I1(\top/processor/sha_core/n586_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10815_12 ),
	.COUT(\top/processor/sha_core/n10814_12 ),
	.SUM(\top/processor/sha_core/n10814_11 )
);
defparam \top/processor/sha_core/n10814_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10813_s3  (
	.I0(\top/processor/sha_core/n10813_7 ),
	.I1(\top/processor/sha_core/n587_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10814_12 ),
	.COUT(\top/processor/sha_core/n10813_12 ),
	.SUM(\top/processor/sha_core/n10813_11 )
);
defparam \top/processor/sha_core/n10813_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10812_s3  (
	.I0(\top/processor/sha_core/n10812_7 ),
	.I1(\top/processor/sha_core/n588_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10813_12 ),
	.COUT(\top/processor/sha_core/n10812_12 ),
	.SUM(\top/processor/sha_core/n10812_11 )
);
defparam \top/processor/sha_core/n10812_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10811_s3  (
	.I0(\top/processor/sha_core/n10811_7 ),
	.I1(\top/processor/sha_core/n589_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10812_12 ),
	.COUT(\top/processor/sha_core/n10811_12 ),
	.SUM(\top/processor/sha_core/n10811_11 )
);
defparam \top/processor/sha_core/n10811_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10810_s3  (
	.I0(\top/processor/sha_core/n10810_7 ),
	.I1(\top/processor/sha_core/n590_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10811_12 ),
	.COUT(\top/processor/sha_core/n10810_12 ),
	.SUM(\top/processor/sha_core/n10810_11 )
);
defparam \top/processor/sha_core/n10810_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10809_s3  (
	.I0(\top/processor/sha_core/n10809_7 ),
	.I1(\top/processor/sha_core/n591_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10810_12 ),
	.COUT(\top/processor/sha_core/n10809_12 ),
	.SUM(\top/processor/sha_core/n10809_11 )
);
defparam \top/processor/sha_core/n10809_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10808_s3  (
	.I0(\top/processor/sha_core/n10808_7 ),
	.I1(\top/processor/sha_core/n592_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10809_12 ),
	.COUT(\top/processor/sha_core/n10808_12 ),
	.SUM(\top/processor/sha_core/n10808_11 )
);
defparam \top/processor/sha_core/n10808_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10807_s3  (
	.I0(\top/processor/sha_core/n10807_7 ),
	.I1(\top/processor/sha_core/n593_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10808_12 ),
	.COUT(\top/processor/sha_core/n10807_12 ),
	.SUM(\top/processor/sha_core/n10807_11 )
);
defparam \top/processor/sha_core/n10807_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10806_s3  (
	.I0(\top/processor/sha_core/n10806_7 ),
	.I1(\top/processor/sha_core/n594_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10807_12 ),
	.COUT(\top/processor/sha_core/n10806_12 ),
	.SUM(\top/processor/sha_core/n10806_11 )
);
defparam \top/processor/sha_core/n10806_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10805_s3  (
	.I0(\top/processor/sha_core/n10805_7 ),
	.I1(\top/processor/sha_core/n595_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10806_12 ),
	.COUT(\top/processor/sha_core/n10805_12 ),
	.SUM(\top/processor/sha_core/n10805_11 )
);
defparam \top/processor/sha_core/n10805_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10804_s3  (
	.I0(\top/processor/sha_core/n10804_7 ),
	.I1(\top/processor/sha_core/n596_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10805_12 ),
	.COUT(\top/processor/sha_core/n10804_12 ),
	.SUM(\top/processor/sha_core/n10804_11 )
);
defparam \top/processor/sha_core/n10804_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10803_s3  (
	.I0(\top/processor/sha_core/n10803_7 ),
	.I1(\top/processor/sha_core/n597_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10804_12 ),
	.COUT(\top/processor/sha_core/n10803_12 ),
	.SUM(\top/processor/sha_core/n10803_11 )
);
defparam \top/processor/sha_core/n10803_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10802_s3  (
	.I0(\top/processor/sha_core/n10802_7 ),
	.I1(\top/processor/sha_core/n598_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10803_12 ),
	.COUT(\top/processor/sha_core/n10802_12 ),
	.SUM(\top/processor/sha_core/n10802_11 )
);
defparam \top/processor/sha_core/n10802_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10801_s3  (
	.I0(\top/processor/sha_core/n10801_7 ),
	.I1(\top/processor/sha_core/n599_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10802_12 ),
	.COUT(\top/processor/sha_core/n10801_12 ),
	.SUM(\top/processor/sha_core/n10801_11 )
);
defparam \top/processor/sha_core/n10801_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10800_s3  (
	.I0(\top/processor/sha_core/n10800_7 ),
	.I1(\top/processor/sha_core/n600_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10801_12 ),
	.COUT(\top/processor/sha_core/n10800_12 ),
	.SUM(\top/processor/sha_core/n10800_11 )
);
defparam \top/processor/sha_core/n10800_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10799_s3  (
	.I0(\top/processor/sha_core/n10799_7 ),
	.I1(\top/processor/sha_core/n601_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10800_12 ),
	.COUT(\top/processor/sha_core/n10799_12 ),
	.SUM(\top/processor/sha_core/n10799_11 )
);
defparam \top/processor/sha_core/n10799_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10798_s3  (
	.I0(\top/processor/sha_core/n10798_7 ),
	.I1(\top/processor/sha_core/n602_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10799_12 ),
	.COUT(\top/processor/sha_core/n10798_12 ),
	.SUM(\top/processor/sha_core/n10798_11 )
);
defparam \top/processor/sha_core/n10798_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10797_s3  (
	.I0(\top/processor/sha_core/n10797_7 ),
	.I1(\top/processor/sha_core/n603_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10798_12 ),
	.COUT(\top/processor/sha_core/n10797_12 ),
	.SUM(\top/processor/sha_core/n10797_11 )
);
defparam \top/processor/sha_core/n10797_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10796_s3  (
	.I0(\top/processor/sha_core/n10796_7 ),
	.I1(\top/processor/sha_core/n604_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10797_12 ),
	.COUT(\top/processor/sha_core/n10796_12 ),
	.SUM(\top/processor/sha_core/n10796_11 )
);
defparam \top/processor/sha_core/n10796_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10795_s3  (
	.I0(\top/processor/sha_core/n10795_7 ),
	.I1(\top/processor/sha_core/n605_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10796_12 ),
	.COUT(\top/processor/sha_core/n10795_12 ),
	.SUM(\top/processor/sha_core/n10795_11 )
);
defparam \top/processor/sha_core/n10795_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10794_s3  (
	.I0(\top/processor/sha_core/n10794_7 ),
	.I1(\top/processor/sha_core/n606_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10795_12 ),
	.COUT(\top/processor/sha_core/n10794_12 ),
	.SUM(\top/processor/sha_core/n10794_11 )
);
defparam \top/processor/sha_core/n10794_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10793_s3  (
	.I0(\top/processor/sha_core/n10793_7 ),
	.I1(\top/processor/sha_core/n607_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10794_12 ),
	.COUT(\top/processor/sha_core/n10793_12 ),
	.SUM(\top/processor/sha_core/n10793_11 )
);
defparam \top/processor/sha_core/n10793_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10792_s3  (
	.I0(\top/processor/sha_core/n10792_7 ),
	.I1(\top/processor/sha_core/n608_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10793_12 ),
	.COUT(\top/processor/sha_core/n10792_12 ),
	.SUM(\top/processor/sha_core/n10792_11 )
);
defparam \top/processor/sha_core/n10792_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10791_s3  (
	.I0(\top/processor/sha_core/n10791_7 ),
	.I1(\top/processor/sha_core/n609_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10792_12 ),
	.COUT(\top/processor/sha_core/n10791_12 ),
	.SUM(\top/processor/sha_core/n10791_11 )
);
defparam \top/processor/sha_core/n10791_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10790_s3  (
	.I0(\top/processor/sha_core/n10790_7 ),
	.I1(\top/processor/sha_core/n610_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10791_12 ),
	.COUT(\top/processor/sha_core/n10790_12 ),
	.SUM(\top/processor/sha_core/n10790_11 )
);
defparam \top/processor/sha_core/n10790_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10789_s3  (
	.I0(\top/processor/sha_core/n10789_7 ),
	.I1(\top/processor/sha_core/n611_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10790_12 ),
	.COUT(\top/processor/sha_core/n10789_12 ),
	.SUM(\top/processor/sha_core/n10789_11 )
);
defparam \top/processor/sha_core/n10789_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10788_s3  (
	.I0(\top/processor/sha_core/n10788_7 ),
	.I1(\top/processor/sha_core/n612_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10789_12 ),
	.COUT(\top/processor/sha_core/n10788_12 ),
	.SUM(\top/processor/sha_core/n10788_11 )
);
defparam \top/processor/sha_core/n10788_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10787_s3  (
	.I0(\top/processor/sha_core/n10787_7 ),
	.I1(\top/processor/sha_core/n613_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10788_12 ),
	.COUT(\top/processor/sha_core/n10787_12 ),
	.SUM(\top/processor/sha_core/n10787_11 )
);
defparam \top/processor/sha_core/n10787_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10786_s3  (
	.I0(\top/processor/sha_core/n10786_7 ),
	.I1(\top/processor/sha_core/n614_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10787_12 ),
	.COUT(\top/processor/sha_core/n10786_12 ),
	.SUM(\top/processor/sha_core/n10786_11 )
);
defparam \top/processor/sha_core/n10786_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10785_s3  (
	.I0(\top/processor/sha_core/n10785_7 ),
	.I1(\top/processor/sha_core/n615_3 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10786_12 ),
	.COUT(\top/processor/sha_core/n10785_4_COUT ),
	.SUM(\top/processor/sha_core/n10785_11 )
);
defparam \top/processor/sha_core/n10785_s3 .ALU_MODE=0;
ALU \top/processor/sha_core/n10816_s4  (
	.I0(\top/processor/sha_core/n10816_9 ),
	.I1(\top/processor/sha_core/n10816_11 ),
	.I3(GND),
	.CIN(GND),
	.COUT(\top/processor/sha_core/n10816_14 ),
	.SUM(\top/processor/sha_core/n10816_13 )
);
defparam \top/processor/sha_core/n10816_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10815_s4  (
	.I0(\top/processor/sha_core/n10815_9 ),
	.I1(\top/processor/sha_core/n10815_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10816_14 ),
	.COUT(\top/processor/sha_core/n10815_14 ),
	.SUM(\top/processor/sha_core/n10815_13 )
);
defparam \top/processor/sha_core/n10815_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10814_s4  (
	.I0(\top/processor/sha_core/n10814_9 ),
	.I1(\top/processor/sha_core/n10814_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10815_14 ),
	.COUT(\top/processor/sha_core/n10814_14 ),
	.SUM(\top/processor/sha_core/n10814_13 )
);
defparam \top/processor/sha_core/n10814_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10813_s4  (
	.I0(\top/processor/sha_core/n10813_9 ),
	.I1(\top/processor/sha_core/n10813_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10814_14 ),
	.COUT(\top/processor/sha_core/n10813_14 ),
	.SUM(\top/processor/sha_core/n10813_13 )
);
defparam \top/processor/sha_core/n10813_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10812_s4  (
	.I0(\top/processor/sha_core/n10812_9 ),
	.I1(\top/processor/sha_core/n10812_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10813_14 ),
	.COUT(\top/processor/sha_core/n10812_14 ),
	.SUM(\top/processor/sha_core/n10812_13 )
);
defparam \top/processor/sha_core/n10812_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10811_s4  (
	.I0(\top/processor/sha_core/n10811_9 ),
	.I1(\top/processor/sha_core/n10811_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10812_14 ),
	.COUT(\top/processor/sha_core/n10811_14 ),
	.SUM(\top/processor/sha_core/n10811_13 )
);
defparam \top/processor/sha_core/n10811_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10810_s4  (
	.I0(\top/processor/sha_core/n10810_9 ),
	.I1(\top/processor/sha_core/n10810_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10811_14 ),
	.COUT(\top/processor/sha_core/n10810_14 ),
	.SUM(\top/processor/sha_core/n10810_13 )
);
defparam \top/processor/sha_core/n10810_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10809_s4  (
	.I0(\top/processor/sha_core/n10809_9 ),
	.I1(\top/processor/sha_core/n10809_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10810_14 ),
	.COUT(\top/processor/sha_core/n10809_14 ),
	.SUM(\top/processor/sha_core/n10809_13 )
);
defparam \top/processor/sha_core/n10809_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10808_s4  (
	.I0(\top/processor/sha_core/n10808_9 ),
	.I1(\top/processor/sha_core/n10808_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10809_14 ),
	.COUT(\top/processor/sha_core/n10808_14 ),
	.SUM(\top/processor/sha_core/n10808_13 )
);
defparam \top/processor/sha_core/n10808_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10807_s4  (
	.I0(\top/processor/sha_core/n10807_9 ),
	.I1(\top/processor/sha_core/n10807_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10808_14 ),
	.COUT(\top/processor/sha_core/n10807_14 ),
	.SUM(\top/processor/sha_core/n10807_13 )
);
defparam \top/processor/sha_core/n10807_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10806_s4  (
	.I0(\top/processor/sha_core/n10806_9 ),
	.I1(\top/processor/sha_core/n10806_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10807_14 ),
	.COUT(\top/processor/sha_core/n10806_14 ),
	.SUM(\top/processor/sha_core/n10806_13 )
);
defparam \top/processor/sha_core/n10806_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10805_s4  (
	.I0(\top/processor/sha_core/n10805_9 ),
	.I1(\top/processor/sha_core/n10805_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10806_14 ),
	.COUT(\top/processor/sha_core/n10805_14 ),
	.SUM(\top/processor/sha_core/n10805_13 )
);
defparam \top/processor/sha_core/n10805_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10804_s4  (
	.I0(\top/processor/sha_core/n10804_9 ),
	.I1(\top/processor/sha_core/n10804_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10805_14 ),
	.COUT(\top/processor/sha_core/n10804_14 ),
	.SUM(\top/processor/sha_core/n10804_13 )
);
defparam \top/processor/sha_core/n10804_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10803_s4  (
	.I0(\top/processor/sha_core/n10803_9 ),
	.I1(\top/processor/sha_core/n10803_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10804_14 ),
	.COUT(\top/processor/sha_core/n10803_14 ),
	.SUM(\top/processor/sha_core/n10803_13 )
);
defparam \top/processor/sha_core/n10803_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10802_s4  (
	.I0(\top/processor/sha_core/n10802_9 ),
	.I1(\top/processor/sha_core/n10802_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10803_14 ),
	.COUT(\top/processor/sha_core/n10802_14 ),
	.SUM(\top/processor/sha_core/n10802_13 )
);
defparam \top/processor/sha_core/n10802_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10801_s4  (
	.I0(\top/processor/sha_core/n10801_9 ),
	.I1(\top/processor/sha_core/n10801_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10802_14 ),
	.COUT(\top/processor/sha_core/n10801_14 ),
	.SUM(\top/processor/sha_core/n10801_13 )
);
defparam \top/processor/sha_core/n10801_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10800_s4  (
	.I0(\top/processor/sha_core/n10800_9 ),
	.I1(\top/processor/sha_core/n10800_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10801_14 ),
	.COUT(\top/processor/sha_core/n10800_14 ),
	.SUM(\top/processor/sha_core/n10800_13 )
);
defparam \top/processor/sha_core/n10800_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10799_s4  (
	.I0(\top/processor/sha_core/n10799_9 ),
	.I1(\top/processor/sha_core/n10799_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10800_14 ),
	.COUT(\top/processor/sha_core/n10799_14 ),
	.SUM(\top/processor/sha_core/n10799_13 )
);
defparam \top/processor/sha_core/n10799_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10798_s4  (
	.I0(\top/processor/sha_core/n10798_9 ),
	.I1(\top/processor/sha_core/n10798_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10799_14 ),
	.COUT(\top/processor/sha_core/n10798_14 ),
	.SUM(\top/processor/sha_core/n10798_13 )
);
defparam \top/processor/sha_core/n10798_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10797_s4  (
	.I0(\top/processor/sha_core/n10797_9 ),
	.I1(\top/processor/sha_core/n10797_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10798_14 ),
	.COUT(\top/processor/sha_core/n10797_14 ),
	.SUM(\top/processor/sha_core/n10797_13 )
);
defparam \top/processor/sha_core/n10797_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10796_s4  (
	.I0(\top/processor/sha_core/n10796_9 ),
	.I1(\top/processor/sha_core/n10796_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10797_14 ),
	.COUT(\top/processor/sha_core/n10796_14 ),
	.SUM(\top/processor/sha_core/n10796_13 )
);
defparam \top/processor/sha_core/n10796_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10795_s4  (
	.I0(\top/processor/sha_core/n10795_9 ),
	.I1(\top/processor/sha_core/n10795_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10796_14 ),
	.COUT(\top/processor/sha_core/n10795_14 ),
	.SUM(\top/processor/sha_core/n10795_13 )
);
defparam \top/processor/sha_core/n10795_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10794_s4  (
	.I0(\top/processor/sha_core/n10794_9 ),
	.I1(\top/processor/sha_core/n10794_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10795_14 ),
	.COUT(\top/processor/sha_core/n10794_14 ),
	.SUM(\top/processor/sha_core/n10794_13 )
);
defparam \top/processor/sha_core/n10794_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10793_s4  (
	.I0(\top/processor/sha_core/n10793_9 ),
	.I1(\top/processor/sha_core/n10793_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10794_14 ),
	.COUT(\top/processor/sha_core/n10793_14 ),
	.SUM(\top/processor/sha_core/n10793_13 )
);
defparam \top/processor/sha_core/n10793_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10792_s4  (
	.I0(\top/processor/sha_core/n10792_9 ),
	.I1(\top/processor/sha_core/n10792_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10793_14 ),
	.COUT(\top/processor/sha_core/n10792_14 ),
	.SUM(\top/processor/sha_core/n10792_13 )
);
defparam \top/processor/sha_core/n10792_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10791_s4  (
	.I0(\top/processor/sha_core/n10791_9 ),
	.I1(\top/processor/sha_core/n10791_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10792_14 ),
	.COUT(\top/processor/sha_core/n10791_14 ),
	.SUM(\top/processor/sha_core/n10791_13 )
);
defparam \top/processor/sha_core/n10791_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10790_s4  (
	.I0(\top/processor/sha_core/n10790_9 ),
	.I1(\top/processor/sha_core/n10790_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10791_14 ),
	.COUT(\top/processor/sha_core/n10790_14 ),
	.SUM(\top/processor/sha_core/n10790_13 )
);
defparam \top/processor/sha_core/n10790_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10789_s4  (
	.I0(\top/processor/sha_core/n10789_9 ),
	.I1(\top/processor/sha_core/n10789_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10790_14 ),
	.COUT(\top/processor/sha_core/n10789_14 ),
	.SUM(\top/processor/sha_core/n10789_13 )
);
defparam \top/processor/sha_core/n10789_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10788_s4  (
	.I0(\top/processor/sha_core/n10788_9 ),
	.I1(\top/processor/sha_core/n10788_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10789_14 ),
	.COUT(\top/processor/sha_core/n10788_14 ),
	.SUM(\top/processor/sha_core/n10788_13 )
);
defparam \top/processor/sha_core/n10788_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10787_s4  (
	.I0(\top/processor/sha_core/n10787_9 ),
	.I1(\top/processor/sha_core/n10787_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10788_14 ),
	.COUT(\top/processor/sha_core/n10787_14 ),
	.SUM(\top/processor/sha_core/n10787_13 )
);
defparam \top/processor/sha_core/n10787_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10786_s4  (
	.I0(\top/processor/sha_core/n10786_9 ),
	.I1(\top/processor/sha_core/n10786_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10787_14 ),
	.COUT(\top/processor/sha_core/n10786_14 ),
	.SUM(\top/processor/sha_core/n10786_13 )
);
defparam \top/processor/sha_core/n10786_s4 .ALU_MODE=0;
ALU \top/processor/sha_core/n10785_s4  (
	.I0(\top/processor/sha_core/n10785_9 ),
	.I1(\top/processor/sha_core/n10785_11 ),
	.I3(GND),
	.CIN(\top/processor/sha_core/n10786_14 ),
	.COUT(\top/processor/sha_core/n10785_5_COUT ),
	.SUM(\top/processor/sha_core/n10785_13 )
);
defparam \top/processor/sha_core/n10785_s4 .ALU_MODE=0;
MUX2_LUT5 \top/processor/sha_core/n327_s202  (
	.I0(\top/processor/sha_core/n327_132 ),
	.I1(\top/processor/sha_core/n327_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_165 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s203  (
	.I0(\top/processor/sha_core/n327_134 ),
	.I1(\top/processor/sha_core/n327_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_167 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s204  (
	.I0(\top/processor/sha_core/n327_136 ),
	.I1(\top/processor/sha_core/n327_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_169 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s205  (
	.I0(\top/processor/sha_core/n327_138 ),
	.I1(\top/processor/sha_core/n327_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_171 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s206  (
	.I0(\top/processor/sha_core/n327_140 ),
	.I1(\top/processor/sha_core/n327_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_173 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s207  (
	.I0(\top/processor/sha_core/n327_142 ),
	.I1(\top/processor/sha_core/n327_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_175 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s208  (
	.I0(\top/processor/sha_core/n327_144 ),
	.I1(\top/processor/sha_core/n327_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_177 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s209  (
	.I0(\top/processor/sha_core/n327_146 ),
	.I1(\top/processor/sha_core/n327_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_179 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s210  (
	.I0(\top/processor/sha_core/n327_148 ),
	.I1(\top/processor/sha_core/n327_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_181 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s211  (
	.I0(\top/processor/sha_core/n327_150 ),
	.I1(\top/processor/sha_core/n327_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_183 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s212  (
	.I0(\top/processor/sha_core/n327_152 ),
	.I1(\top/processor/sha_core/n327_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_185 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s213  (
	.I0(\top/processor/sha_core/n327_154 ),
	.I1(\top/processor/sha_core/n327_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_187 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s214  (
	.I0(\top/processor/sha_core/n327_156 ),
	.I1(\top/processor/sha_core/n327_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_189 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s215  (
	.I0(\top/processor/sha_core/n327_158 ),
	.I1(\top/processor/sha_core/n327_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_191 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s216  (
	.I0(\top/processor/sha_core/n327_160 ),
	.I1(\top/processor/sha_core/n327_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_193 )
);
MUX2_LUT5 \top/processor/sha_core/n327_s217  (
	.I0(\top/processor/sha_core/n327_162 ),
	.I1(\top/processor/sha_core/n327_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n327_195 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s202  (
	.I0(\top/processor/sha_core/n328_132 ),
	.I1(\top/processor/sha_core/n328_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_165 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s203  (
	.I0(\top/processor/sha_core/n328_134 ),
	.I1(\top/processor/sha_core/n328_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_167 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s204  (
	.I0(\top/processor/sha_core/n328_136 ),
	.I1(\top/processor/sha_core/n328_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_169 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s205  (
	.I0(\top/processor/sha_core/n328_138 ),
	.I1(\top/processor/sha_core/n328_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_171 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s206  (
	.I0(\top/processor/sha_core/n328_140 ),
	.I1(\top/processor/sha_core/n328_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_173 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s207  (
	.I0(\top/processor/sha_core/n328_142 ),
	.I1(\top/processor/sha_core/n328_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_175 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s208  (
	.I0(\top/processor/sha_core/n328_144 ),
	.I1(\top/processor/sha_core/n328_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_177 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s209  (
	.I0(\top/processor/sha_core/n328_146 ),
	.I1(\top/processor/sha_core/n328_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_179 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s210  (
	.I0(\top/processor/sha_core/n328_148 ),
	.I1(\top/processor/sha_core/n328_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_181 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s211  (
	.I0(\top/processor/sha_core/n328_150 ),
	.I1(\top/processor/sha_core/n328_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_183 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s212  (
	.I0(\top/processor/sha_core/n328_152 ),
	.I1(\top/processor/sha_core/n328_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_185 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s213  (
	.I0(\top/processor/sha_core/n328_154 ),
	.I1(\top/processor/sha_core/n328_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_187 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s214  (
	.I0(\top/processor/sha_core/n328_156 ),
	.I1(\top/processor/sha_core/n328_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_189 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s215  (
	.I0(\top/processor/sha_core/n328_158 ),
	.I1(\top/processor/sha_core/n328_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_191 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s216  (
	.I0(\top/processor/sha_core/n328_160 ),
	.I1(\top/processor/sha_core/n328_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_193 )
);
MUX2_LUT5 \top/processor/sha_core/n328_s217  (
	.I0(\top/processor/sha_core/n328_162 ),
	.I1(\top/processor/sha_core/n328_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n328_195 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s202  (
	.I0(\top/processor/sha_core/n329_132 ),
	.I1(\top/processor/sha_core/n329_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_165 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s203  (
	.I0(\top/processor/sha_core/n329_134 ),
	.I1(\top/processor/sha_core/n329_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_167 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s204  (
	.I0(\top/processor/sha_core/n329_136 ),
	.I1(\top/processor/sha_core/n329_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_169 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s205  (
	.I0(\top/processor/sha_core/n329_138 ),
	.I1(\top/processor/sha_core/n329_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_171 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s206  (
	.I0(\top/processor/sha_core/n329_140 ),
	.I1(\top/processor/sha_core/n329_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_173 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s207  (
	.I0(\top/processor/sha_core/n329_142 ),
	.I1(\top/processor/sha_core/n329_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_175 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s208  (
	.I0(\top/processor/sha_core/n329_144 ),
	.I1(\top/processor/sha_core/n329_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_177 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s209  (
	.I0(\top/processor/sha_core/n329_146 ),
	.I1(\top/processor/sha_core/n329_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_179 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s210  (
	.I0(\top/processor/sha_core/n329_148 ),
	.I1(\top/processor/sha_core/n329_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_181 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s211  (
	.I0(\top/processor/sha_core/n329_150 ),
	.I1(\top/processor/sha_core/n329_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_183 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s212  (
	.I0(\top/processor/sha_core/n329_152 ),
	.I1(\top/processor/sha_core/n329_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_185 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s213  (
	.I0(\top/processor/sha_core/n329_154 ),
	.I1(\top/processor/sha_core/n329_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_187 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s214  (
	.I0(\top/processor/sha_core/n329_156 ),
	.I1(\top/processor/sha_core/n329_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_189 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s215  (
	.I0(\top/processor/sha_core/n329_158 ),
	.I1(\top/processor/sha_core/n329_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_191 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s216  (
	.I0(\top/processor/sha_core/n329_160 ),
	.I1(\top/processor/sha_core/n329_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_193 )
);
MUX2_LUT5 \top/processor/sha_core/n329_s217  (
	.I0(\top/processor/sha_core/n329_162 ),
	.I1(\top/processor/sha_core/n329_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n329_195 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s202  (
	.I0(\top/processor/sha_core/n330_132 ),
	.I1(\top/processor/sha_core/n330_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_165 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s203  (
	.I0(\top/processor/sha_core/n330_134 ),
	.I1(\top/processor/sha_core/n330_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_167 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s204  (
	.I0(\top/processor/sha_core/n330_136 ),
	.I1(\top/processor/sha_core/n330_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_169 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s205  (
	.I0(\top/processor/sha_core/n330_138 ),
	.I1(\top/processor/sha_core/n330_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_171 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s206  (
	.I0(\top/processor/sha_core/n330_140 ),
	.I1(\top/processor/sha_core/n330_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_173 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s207  (
	.I0(\top/processor/sha_core/n330_142 ),
	.I1(\top/processor/sha_core/n330_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_175 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s208  (
	.I0(\top/processor/sha_core/n330_144 ),
	.I1(\top/processor/sha_core/n330_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_177 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s209  (
	.I0(\top/processor/sha_core/n330_146 ),
	.I1(\top/processor/sha_core/n330_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_179 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s210  (
	.I0(\top/processor/sha_core/n330_148 ),
	.I1(\top/processor/sha_core/n330_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_181 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s211  (
	.I0(\top/processor/sha_core/n330_150 ),
	.I1(\top/processor/sha_core/n330_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_183 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s212  (
	.I0(\top/processor/sha_core/n330_152 ),
	.I1(\top/processor/sha_core/n330_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_185 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s213  (
	.I0(\top/processor/sha_core/n330_154 ),
	.I1(\top/processor/sha_core/n330_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_187 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s214  (
	.I0(\top/processor/sha_core/n330_156 ),
	.I1(\top/processor/sha_core/n330_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_189 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s215  (
	.I0(\top/processor/sha_core/n330_158 ),
	.I1(\top/processor/sha_core/n330_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_191 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s216  (
	.I0(\top/processor/sha_core/n330_160 ),
	.I1(\top/processor/sha_core/n330_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_193 )
);
MUX2_LUT5 \top/processor/sha_core/n330_s217  (
	.I0(\top/processor/sha_core/n330_162 ),
	.I1(\top/processor/sha_core/n330_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n330_195 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s202  (
	.I0(\top/processor/sha_core/n331_132 ),
	.I1(\top/processor/sha_core/n331_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_165 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s203  (
	.I0(\top/processor/sha_core/n331_134 ),
	.I1(\top/processor/sha_core/n331_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_167 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s204  (
	.I0(\top/processor/sha_core/n331_136 ),
	.I1(\top/processor/sha_core/n331_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_169 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s205  (
	.I0(\top/processor/sha_core/n331_138 ),
	.I1(\top/processor/sha_core/n331_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_171 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s206  (
	.I0(\top/processor/sha_core/n331_140 ),
	.I1(\top/processor/sha_core/n331_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_173 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s207  (
	.I0(\top/processor/sha_core/n331_142 ),
	.I1(\top/processor/sha_core/n331_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_175 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s208  (
	.I0(\top/processor/sha_core/n331_144 ),
	.I1(\top/processor/sha_core/n331_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_177 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s209  (
	.I0(\top/processor/sha_core/n331_146 ),
	.I1(\top/processor/sha_core/n331_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_179 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s210  (
	.I0(\top/processor/sha_core/n331_148 ),
	.I1(\top/processor/sha_core/n331_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_181 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s211  (
	.I0(\top/processor/sha_core/n331_150 ),
	.I1(\top/processor/sha_core/n331_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_183 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s212  (
	.I0(\top/processor/sha_core/n331_152 ),
	.I1(\top/processor/sha_core/n331_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_185 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s213  (
	.I0(\top/processor/sha_core/n331_154 ),
	.I1(\top/processor/sha_core/n331_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_187 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s214  (
	.I0(\top/processor/sha_core/n331_156 ),
	.I1(\top/processor/sha_core/n331_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_189 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s215  (
	.I0(\top/processor/sha_core/n331_158 ),
	.I1(\top/processor/sha_core/n331_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_191 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s216  (
	.I0(\top/processor/sha_core/n331_160 ),
	.I1(\top/processor/sha_core/n331_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_193 )
);
MUX2_LUT5 \top/processor/sha_core/n331_s217  (
	.I0(\top/processor/sha_core/n331_162 ),
	.I1(\top/processor/sha_core/n331_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n331_195 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s202  (
	.I0(\top/processor/sha_core/n332_132 ),
	.I1(\top/processor/sha_core/n332_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_165 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s203  (
	.I0(\top/processor/sha_core/n332_134 ),
	.I1(\top/processor/sha_core/n332_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_167 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s204  (
	.I0(\top/processor/sha_core/n332_136 ),
	.I1(\top/processor/sha_core/n332_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_169 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s205  (
	.I0(\top/processor/sha_core/n332_138 ),
	.I1(\top/processor/sha_core/n332_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_171 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s206  (
	.I0(\top/processor/sha_core/n332_140 ),
	.I1(\top/processor/sha_core/n332_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_173 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s207  (
	.I0(\top/processor/sha_core/n332_142 ),
	.I1(\top/processor/sha_core/n332_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_175 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s208  (
	.I0(\top/processor/sha_core/n332_144 ),
	.I1(\top/processor/sha_core/n332_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_177 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s209  (
	.I0(\top/processor/sha_core/n332_146 ),
	.I1(\top/processor/sha_core/n332_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_179 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s210  (
	.I0(\top/processor/sha_core/n332_148 ),
	.I1(\top/processor/sha_core/n332_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_181 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s211  (
	.I0(\top/processor/sha_core/n332_150 ),
	.I1(\top/processor/sha_core/n332_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_183 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s212  (
	.I0(\top/processor/sha_core/n332_152 ),
	.I1(\top/processor/sha_core/n332_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_185 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s213  (
	.I0(\top/processor/sha_core/n332_154 ),
	.I1(\top/processor/sha_core/n332_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_187 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s214  (
	.I0(\top/processor/sha_core/n332_156 ),
	.I1(\top/processor/sha_core/n332_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_189 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s215  (
	.I0(\top/processor/sha_core/n332_158 ),
	.I1(\top/processor/sha_core/n332_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_191 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s216  (
	.I0(\top/processor/sha_core/n332_160 ),
	.I1(\top/processor/sha_core/n332_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_193 )
);
MUX2_LUT5 \top/processor/sha_core/n332_s217  (
	.I0(\top/processor/sha_core/n332_162 ),
	.I1(\top/processor/sha_core/n332_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n332_195 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s202  (
	.I0(\top/processor/sha_core/n333_132 ),
	.I1(\top/processor/sha_core/n333_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_165 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s203  (
	.I0(\top/processor/sha_core/n333_134 ),
	.I1(\top/processor/sha_core/n333_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_167 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s204  (
	.I0(\top/processor/sha_core/n333_136 ),
	.I1(\top/processor/sha_core/n333_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_169 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s205  (
	.I0(\top/processor/sha_core/n333_138 ),
	.I1(\top/processor/sha_core/n333_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_171 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s206  (
	.I0(\top/processor/sha_core/n333_140 ),
	.I1(\top/processor/sha_core/n333_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_173 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s207  (
	.I0(\top/processor/sha_core/n333_142 ),
	.I1(\top/processor/sha_core/n333_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_175 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s208  (
	.I0(\top/processor/sha_core/n333_144 ),
	.I1(\top/processor/sha_core/n333_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_177 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s209  (
	.I0(\top/processor/sha_core/n333_146 ),
	.I1(\top/processor/sha_core/n333_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_179 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s210  (
	.I0(\top/processor/sha_core/n333_148 ),
	.I1(\top/processor/sha_core/n333_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_181 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s211  (
	.I0(\top/processor/sha_core/n333_150 ),
	.I1(\top/processor/sha_core/n333_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_183 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s212  (
	.I0(\top/processor/sha_core/n333_152 ),
	.I1(\top/processor/sha_core/n333_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_185 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s213  (
	.I0(\top/processor/sha_core/n333_154 ),
	.I1(\top/processor/sha_core/n333_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_187 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s214  (
	.I0(\top/processor/sha_core/n333_156 ),
	.I1(\top/processor/sha_core/n333_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_189 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s215  (
	.I0(\top/processor/sha_core/n333_158 ),
	.I1(\top/processor/sha_core/n333_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_191 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s216  (
	.I0(\top/processor/sha_core/n333_160 ),
	.I1(\top/processor/sha_core/n333_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_193 )
);
MUX2_LUT5 \top/processor/sha_core/n333_s217  (
	.I0(\top/processor/sha_core/n333_162 ),
	.I1(\top/processor/sha_core/n333_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n333_195 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s202  (
	.I0(\top/processor/sha_core/n334_132 ),
	.I1(\top/processor/sha_core/n334_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_165 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s203  (
	.I0(\top/processor/sha_core/n334_134 ),
	.I1(\top/processor/sha_core/n334_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_167 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s204  (
	.I0(\top/processor/sha_core/n334_136 ),
	.I1(\top/processor/sha_core/n334_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_169 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s205  (
	.I0(\top/processor/sha_core/n334_138 ),
	.I1(\top/processor/sha_core/n334_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_171 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s206  (
	.I0(\top/processor/sha_core/n334_140 ),
	.I1(\top/processor/sha_core/n334_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_173 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s207  (
	.I0(\top/processor/sha_core/n334_142 ),
	.I1(\top/processor/sha_core/n334_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_175 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s208  (
	.I0(\top/processor/sha_core/n334_144 ),
	.I1(\top/processor/sha_core/n334_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_177 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s209  (
	.I0(\top/processor/sha_core/n334_146 ),
	.I1(\top/processor/sha_core/n334_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_179 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s210  (
	.I0(\top/processor/sha_core/n334_148 ),
	.I1(\top/processor/sha_core/n334_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_181 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s211  (
	.I0(\top/processor/sha_core/n334_150 ),
	.I1(\top/processor/sha_core/n334_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_183 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s212  (
	.I0(\top/processor/sha_core/n334_152 ),
	.I1(\top/processor/sha_core/n334_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_185 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s213  (
	.I0(\top/processor/sha_core/n334_154 ),
	.I1(\top/processor/sha_core/n334_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_187 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s214  (
	.I0(\top/processor/sha_core/n334_156 ),
	.I1(\top/processor/sha_core/n334_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_189 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s215  (
	.I0(\top/processor/sha_core/n334_158 ),
	.I1(\top/processor/sha_core/n334_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_191 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s216  (
	.I0(\top/processor/sha_core/n334_160 ),
	.I1(\top/processor/sha_core/n334_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_193 )
);
MUX2_LUT5 \top/processor/sha_core/n334_s217  (
	.I0(\top/processor/sha_core/n334_162 ),
	.I1(\top/processor/sha_core/n334_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n334_195 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s202  (
	.I0(\top/processor/sha_core/n335_132 ),
	.I1(\top/processor/sha_core/n335_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_165 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s203  (
	.I0(\top/processor/sha_core/n335_134 ),
	.I1(\top/processor/sha_core/n335_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_167 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s204  (
	.I0(\top/processor/sha_core/n335_136 ),
	.I1(\top/processor/sha_core/n335_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_169 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s205  (
	.I0(\top/processor/sha_core/n335_138 ),
	.I1(\top/processor/sha_core/n335_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_171 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s206  (
	.I0(\top/processor/sha_core/n335_140 ),
	.I1(\top/processor/sha_core/n335_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_173 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s207  (
	.I0(\top/processor/sha_core/n335_142 ),
	.I1(\top/processor/sha_core/n335_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_175 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s208  (
	.I0(\top/processor/sha_core/n335_144 ),
	.I1(\top/processor/sha_core/n335_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_177 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s209  (
	.I0(\top/processor/sha_core/n335_146 ),
	.I1(\top/processor/sha_core/n335_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_179 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s210  (
	.I0(\top/processor/sha_core/n335_148 ),
	.I1(\top/processor/sha_core/n335_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_181 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s211  (
	.I0(\top/processor/sha_core/n335_150 ),
	.I1(\top/processor/sha_core/n335_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_183 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s212  (
	.I0(\top/processor/sha_core/n335_152 ),
	.I1(\top/processor/sha_core/n335_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_185 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s213  (
	.I0(\top/processor/sha_core/n335_154 ),
	.I1(\top/processor/sha_core/n335_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_187 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s214  (
	.I0(\top/processor/sha_core/n335_156 ),
	.I1(\top/processor/sha_core/n335_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_189 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s215  (
	.I0(\top/processor/sha_core/n335_158 ),
	.I1(\top/processor/sha_core/n335_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_191 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s216  (
	.I0(\top/processor/sha_core/n335_160 ),
	.I1(\top/processor/sha_core/n335_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_193 )
);
MUX2_LUT5 \top/processor/sha_core/n335_s217  (
	.I0(\top/processor/sha_core/n335_162 ),
	.I1(\top/processor/sha_core/n335_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n335_195 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s202  (
	.I0(\top/processor/sha_core/n336_132 ),
	.I1(\top/processor/sha_core/n336_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_165 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s203  (
	.I0(\top/processor/sha_core/n336_134 ),
	.I1(\top/processor/sha_core/n336_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_167 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s204  (
	.I0(\top/processor/sha_core/n336_136 ),
	.I1(\top/processor/sha_core/n336_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_169 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s205  (
	.I0(\top/processor/sha_core/n336_138 ),
	.I1(\top/processor/sha_core/n336_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_171 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s206  (
	.I0(\top/processor/sha_core/n336_140 ),
	.I1(\top/processor/sha_core/n336_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_173 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s207  (
	.I0(\top/processor/sha_core/n336_142 ),
	.I1(\top/processor/sha_core/n336_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_175 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s208  (
	.I0(\top/processor/sha_core/n336_144 ),
	.I1(\top/processor/sha_core/n336_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_177 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s209  (
	.I0(\top/processor/sha_core/n336_146 ),
	.I1(\top/processor/sha_core/n336_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_179 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s210  (
	.I0(\top/processor/sha_core/n336_148 ),
	.I1(\top/processor/sha_core/n336_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_181 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s211  (
	.I0(\top/processor/sha_core/n336_150 ),
	.I1(\top/processor/sha_core/n336_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_183 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s212  (
	.I0(\top/processor/sha_core/n336_152 ),
	.I1(\top/processor/sha_core/n336_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_185 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s213  (
	.I0(\top/processor/sha_core/n336_154 ),
	.I1(\top/processor/sha_core/n336_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_187 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s214  (
	.I0(\top/processor/sha_core/n336_156 ),
	.I1(\top/processor/sha_core/n336_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_189 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s215  (
	.I0(\top/processor/sha_core/n336_158 ),
	.I1(\top/processor/sha_core/n336_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_191 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s216  (
	.I0(\top/processor/sha_core/n336_160 ),
	.I1(\top/processor/sha_core/n336_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_193 )
);
MUX2_LUT5 \top/processor/sha_core/n336_s217  (
	.I0(\top/processor/sha_core/n336_162 ),
	.I1(\top/processor/sha_core/n336_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n336_195 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s202  (
	.I0(\top/processor/sha_core/n337_132 ),
	.I1(\top/processor/sha_core/n337_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_165 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s203  (
	.I0(\top/processor/sha_core/n337_134 ),
	.I1(\top/processor/sha_core/n337_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_167 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s204  (
	.I0(\top/processor/sha_core/n337_136 ),
	.I1(\top/processor/sha_core/n337_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_169 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s205  (
	.I0(\top/processor/sha_core/n337_138 ),
	.I1(\top/processor/sha_core/n337_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_171 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s206  (
	.I0(\top/processor/sha_core/n337_140 ),
	.I1(\top/processor/sha_core/n337_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_173 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s207  (
	.I0(\top/processor/sha_core/n337_142 ),
	.I1(\top/processor/sha_core/n337_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_175 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s208  (
	.I0(\top/processor/sha_core/n337_144 ),
	.I1(\top/processor/sha_core/n337_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_177 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s209  (
	.I0(\top/processor/sha_core/n337_146 ),
	.I1(\top/processor/sha_core/n337_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_179 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s210  (
	.I0(\top/processor/sha_core/n337_148 ),
	.I1(\top/processor/sha_core/n337_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_181 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s211  (
	.I0(\top/processor/sha_core/n337_150 ),
	.I1(\top/processor/sha_core/n337_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_183 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s212  (
	.I0(\top/processor/sha_core/n337_152 ),
	.I1(\top/processor/sha_core/n337_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_185 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s213  (
	.I0(\top/processor/sha_core/n337_154 ),
	.I1(\top/processor/sha_core/n337_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_187 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s214  (
	.I0(\top/processor/sha_core/n337_156 ),
	.I1(\top/processor/sha_core/n337_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_189 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s215  (
	.I0(\top/processor/sha_core/n337_158 ),
	.I1(\top/processor/sha_core/n337_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_191 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s216  (
	.I0(\top/processor/sha_core/n337_160 ),
	.I1(\top/processor/sha_core/n337_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_193 )
);
MUX2_LUT5 \top/processor/sha_core/n337_s217  (
	.I0(\top/processor/sha_core/n337_162 ),
	.I1(\top/processor/sha_core/n337_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n337_195 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s202  (
	.I0(\top/processor/sha_core/n338_132 ),
	.I1(\top/processor/sha_core/n338_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_165 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s203  (
	.I0(\top/processor/sha_core/n338_134 ),
	.I1(\top/processor/sha_core/n338_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_167 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s204  (
	.I0(\top/processor/sha_core/n338_136 ),
	.I1(\top/processor/sha_core/n338_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_169 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s205  (
	.I0(\top/processor/sha_core/n338_138 ),
	.I1(\top/processor/sha_core/n338_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_171 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s206  (
	.I0(\top/processor/sha_core/n338_140 ),
	.I1(\top/processor/sha_core/n338_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_173 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s207  (
	.I0(\top/processor/sha_core/n338_142 ),
	.I1(\top/processor/sha_core/n338_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_175 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s208  (
	.I0(\top/processor/sha_core/n338_144 ),
	.I1(\top/processor/sha_core/n338_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_177 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s209  (
	.I0(\top/processor/sha_core/n338_146 ),
	.I1(\top/processor/sha_core/n338_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_179 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s210  (
	.I0(\top/processor/sha_core/n338_148 ),
	.I1(\top/processor/sha_core/n338_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_181 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s211  (
	.I0(\top/processor/sha_core/n338_150 ),
	.I1(\top/processor/sha_core/n338_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_183 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s212  (
	.I0(\top/processor/sha_core/n338_152 ),
	.I1(\top/processor/sha_core/n338_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_185 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s213  (
	.I0(\top/processor/sha_core/n338_154 ),
	.I1(\top/processor/sha_core/n338_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_187 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s214  (
	.I0(\top/processor/sha_core/n338_156 ),
	.I1(\top/processor/sha_core/n338_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_189 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s215  (
	.I0(\top/processor/sha_core/n338_158 ),
	.I1(\top/processor/sha_core/n338_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_191 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s216  (
	.I0(\top/processor/sha_core/n338_160 ),
	.I1(\top/processor/sha_core/n338_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_193 )
);
MUX2_LUT5 \top/processor/sha_core/n338_s217  (
	.I0(\top/processor/sha_core/n338_162 ),
	.I1(\top/processor/sha_core/n338_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n338_195 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s202  (
	.I0(\top/processor/sha_core/n339_132 ),
	.I1(\top/processor/sha_core/n339_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_165 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s203  (
	.I0(\top/processor/sha_core/n339_134 ),
	.I1(\top/processor/sha_core/n339_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_167 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s204  (
	.I0(\top/processor/sha_core/n339_136 ),
	.I1(\top/processor/sha_core/n339_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_169 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s205  (
	.I0(\top/processor/sha_core/n339_138 ),
	.I1(\top/processor/sha_core/n339_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_171 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s206  (
	.I0(\top/processor/sha_core/n339_140 ),
	.I1(\top/processor/sha_core/n339_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_173 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s207  (
	.I0(\top/processor/sha_core/n339_142 ),
	.I1(\top/processor/sha_core/n339_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_175 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s208  (
	.I0(\top/processor/sha_core/n339_144 ),
	.I1(\top/processor/sha_core/n339_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_177 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s209  (
	.I0(\top/processor/sha_core/n339_146 ),
	.I1(\top/processor/sha_core/n339_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_179 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s210  (
	.I0(\top/processor/sha_core/n339_148 ),
	.I1(\top/processor/sha_core/n339_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_181 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s211  (
	.I0(\top/processor/sha_core/n339_150 ),
	.I1(\top/processor/sha_core/n339_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_183 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s212  (
	.I0(\top/processor/sha_core/n339_152 ),
	.I1(\top/processor/sha_core/n339_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_185 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s213  (
	.I0(\top/processor/sha_core/n339_154 ),
	.I1(\top/processor/sha_core/n339_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_187 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s214  (
	.I0(\top/processor/sha_core/n339_156 ),
	.I1(\top/processor/sha_core/n339_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_189 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s215  (
	.I0(\top/processor/sha_core/n339_158 ),
	.I1(\top/processor/sha_core/n339_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_191 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s216  (
	.I0(\top/processor/sha_core/n339_160 ),
	.I1(\top/processor/sha_core/n339_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_193 )
);
MUX2_LUT5 \top/processor/sha_core/n339_s217  (
	.I0(\top/processor/sha_core/n339_162 ),
	.I1(\top/processor/sha_core/n339_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n339_195 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s202  (
	.I0(\top/processor/sha_core/n340_132 ),
	.I1(\top/processor/sha_core/n340_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_165 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s203  (
	.I0(\top/processor/sha_core/n340_134 ),
	.I1(\top/processor/sha_core/n340_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_167 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s204  (
	.I0(\top/processor/sha_core/n340_136 ),
	.I1(\top/processor/sha_core/n340_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_169 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s205  (
	.I0(\top/processor/sha_core/n340_138 ),
	.I1(\top/processor/sha_core/n340_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_171 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s206  (
	.I0(\top/processor/sha_core/n340_140 ),
	.I1(\top/processor/sha_core/n340_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_173 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s207  (
	.I0(\top/processor/sha_core/n340_142 ),
	.I1(\top/processor/sha_core/n340_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_175 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s208  (
	.I0(\top/processor/sha_core/n340_144 ),
	.I1(\top/processor/sha_core/n340_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_177 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s209  (
	.I0(\top/processor/sha_core/n340_146 ),
	.I1(\top/processor/sha_core/n340_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_179 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s210  (
	.I0(\top/processor/sha_core/n340_148 ),
	.I1(\top/processor/sha_core/n340_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_181 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s211  (
	.I0(\top/processor/sha_core/n340_150 ),
	.I1(\top/processor/sha_core/n340_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_183 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s212  (
	.I0(\top/processor/sha_core/n340_152 ),
	.I1(\top/processor/sha_core/n340_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_185 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s213  (
	.I0(\top/processor/sha_core/n340_154 ),
	.I1(\top/processor/sha_core/n340_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_187 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s214  (
	.I0(\top/processor/sha_core/n340_156 ),
	.I1(\top/processor/sha_core/n340_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_189 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s215  (
	.I0(\top/processor/sha_core/n340_158 ),
	.I1(\top/processor/sha_core/n340_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_191 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s216  (
	.I0(\top/processor/sha_core/n340_160 ),
	.I1(\top/processor/sha_core/n340_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_193 )
);
MUX2_LUT5 \top/processor/sha_core/n340_s217  (
	.I0(\top/processor/sha_core/n340_162 ),
	.I1(\top/processor/sha_core/n340_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n340_195 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s202  (
	.I0(\top/processor/sha_core/n341_132 ),
	.I1(\top/processor/sha_core/n341_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_165 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s203  (
	.I0(\top/processor/sha_core/n341_134 ),
	.I1(\top/processor/sha_core/n341_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_167 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s204  (
	.I0(\top/processor/sha_core/n341_136 ),
	.I1(\top/processor/sha_core/n341_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_169 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s205  (
	.I0(\top/processor/sha_core/n341_138 ),
	.I1(\top/processor/sha_core/n341_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_171 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s206  (
	.I0(\top/processor/sha_core/n341_140 ),
	.I1(\top/processor/sha_core/n341_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_173 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s207  (
	.I0(\top/processor/sha_core/n341_142 ),
	.I1(\top/processor/sha_core/n341_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_175 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s208  (
	.I0(\top/processor/sha_core/n341_144 ),
	.I1(\top/processor/sha_core/n341_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_177 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s209  (
	.I0(\top/processor/sha_core/n341_146 ),
	.I1(\top/processor/sha_core/n341_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_179 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s210  (
	.I0(\top/processor/sha_core/n341_148 ),
	.I1(\top/processor/sha_core/n341_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_181 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s211  (
	.I0(\top/processor/sha_core/n341_150 ),
	.I1(\top/processor/sha_core/n341_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_183 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s212  (
	.I0(\top/processor/sha_core/n341_152 ),
	.I1(\top/processor/sha_core/n341_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_185 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s213  (
	.I0(\top/processor/sha_core/n341_154 ),
	.I1(\top/processor/sha_core/n341_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_187 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s214  (
	.I0(\top/processor/sha_core/n341_156 ),
	.I1(\top/processor/sha_core/n341_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_189 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s215  (
	.I0(\top/processor/sha_core/n341_158 ),
	.I1(\top/processor/sha_core/n341_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_191 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s216  (
	.I0(\top/processor/sha_core/n341_160 ),
	.I1(\top/processor/sha_core/n341_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_193 )
);
MUX2_LUT5 \top/processor/sha_core/n341_s217  (
	.I0(\top/processor/sha_core/n341_162 ),
	.I1(\top/processor/sha_core/n341_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n341_195 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s202  (
	.I0(\top/processor/sha_core/n342_132 ),
	.I1(\top/processor/sha_core/n342_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_165 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s203  (
	.I0(\top/processor/sha_core/n342_134 ),
	.I1(\top/processor/sha_core/n342_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_167 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s204  (
	.I0(\top/processor/sha_core/n342_136 ),
	.I1(\top/processor/sha_core/n342_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_169 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s205  (
	.I0(\top/processor/sha_core/n342_138 ),
	.I1(\top/processor/sha_core/n342_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_171 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s206  (
	.I0(\top/processor/sha_core/n342_140 ),
	.I1(\top/processor/sha_core/n342_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_173 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s207  (
	.I0(\top/processor/sha_core/n342_142 ),
	.I1(\top/processor/sha_core/n342_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_175 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s208  (
	.I0(\top/processor/sha_core/n342_144 ),
	.I1(\top/processor/sha_core/n342_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_177 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s209  (
	.I0(\top/processor/sha_core/n342_146 ),
	.I1(\top/processor/sha_core/n342_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_179 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s210  (
	.I0(\top/processor/sha_core/n342_148 ),
	.I1(\top/processor/sha_core/n342_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_181 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s211  (
	.I0(\top/processor/sha_core/n342_150 ),
	.I1(\top/processor/sha_core/n342_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_183 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s212  (
	.I0(\top/processor/sha_core/n342_152 ),
	.I1(\top/processor/sha_core/n342_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_185 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s213  (
	.I0(\top/processor/sha_core/n342_154 ),
	.I1(\top/processor/sha_core/n342_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_187 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s214  (
	.I0(\top/processor/sha_core/n342_156 ),
	.I1(\top/processor/sha_core/n342_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_189 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s215  (
	.I0(\top/processor/sha_core/n342_158 ),
	.I1(\top/processor/sha_core/n342_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_191 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s216  (
	.I0(\top/processor/sha_core/n342_160 ),
	.I1(\top/processor/sha_core/n342_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_193 )
);
MUX2_LUT5 \top/processor/sha_core/n342_s217  (
	.I0(\top/processor/sha_core/n342_162 ),
	.I1(\top/processor/sha_core/n342_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n342_195 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s202  (
	.I0(\top/processor/sha_core/n343_132 ),
	.I1(\top/processor/sha_core/n343_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_165 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s203  (
	.I0(\top/processor/sha_core/n343_134 ),
	.I1(\top/processor/sha_core/n343_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_167 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s204  (
	.I0(\top/processor/sha_core/n343_136 ),
	.I1(\top/processor/sha_core/n343_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_169 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s205  (
	.I0(\top/processor/sha_core/n343_138 ),
	.I1(\top/processor/sha_core/n343_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_171 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s206  (
	.I0(\top/processor/sha_core/n343_140 ),
	.I1(\top/processor/sha_core/n343_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_173 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s207  (
	.I0(\top/processor/sha_core/n343_142 ),
	.I1(\top/processor/sha_core/n343_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_175 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s208  (
	.I0(\top/processor/sha_core/n343_144 ),
	.I1(\top/processor/sha_core/n343_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_177 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s209  (
	.I0(\top/processor/sha_core/n343_146 ),
	.I1(\top/processor/sha_core/n343_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_179 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s210  (
	.I0(\top/processor/sha_core/n343_148 ),
	.I1(\top/processor/sha_core/n343_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_181 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s211  (
	.I0(\top/processor/sha_core/n343_150 ),
	.I1(\top/processor/sha_core/n343_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_183 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s212  (
	.I0(\top/processor/sha_core/n343_152 ),
	.I1(\top/processor/sha_core/n343_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_185 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s213  (
	.I0(\top/processor/sha_core/n343_154 ),
	.I1(\top/processor/sha_core/n343_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_187 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s214  (
	.I0(\top/processor/sha_core/n343_156 ),
	.I1(\top/processor/sha_core/n343_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_189 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s215  (
	.I0(\top/processor/sha_core/n343_158 ),
	.I1(\top/processor/sha_core/n343_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_191 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s216  (
	.I0(\top/processor/sha_core/n343_160 ),
	.I1(\top/processor/sha_core/n343_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_193 )
);
MUX2_LUT5 \top/processor/sha_core/n343_s217  (
	.I0(\top/processor/sha_core/n343_162 ),
	.I1(\top/processor/sha_core/n343_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n343_195 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s202  (
	.I0(\top/processor/sha_core/n344_132 ),
	.I1(\top/processor/sha_core/n344_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_165 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s203  (
	.I0(\top/processor/sha_core/n344_134 ),
	.I1(\top/processor/sha_core/n344_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_167 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s204  (
	.I0(\top/processor/sha_core/n344_136 ),
	.I1(\top/processor/sha_core/n344_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_169 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s205  (
	.I0(\top/processor/sha_core/n344_138 ),
	.I1(\top/processor/sha_core/n344_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_171 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s206  (
	.I0(\top/processor/sha_core/n344_140 ),
	.I1(\top/processor/sha_core/n344_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_173 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s207  (
	.I0(\top/processor/sha_core/n344_142 ),
	.I1(\top/processor/sha_core/n344_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_175 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s208  (
	.I0(\top/processor/sha_core/n344_144 ),
	.I1(\top/processor/sha_core/n344_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_177 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s209  (
	.I0(\top/processor/sha_core/n344_146 ),
	.I1(\top/processor/sha_core/n344_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_179 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s210  (
	.I0(\top/processor/sha_core/n344_148 ),
	.I1(\top/processor/sha_core/n344_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_181 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s211  (
	.I0(\top/processor/sha_core/n344_150 ),
	.I1(\top/processor/sha_core/n344_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_183 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s212  (
	.I0(\top/processor/sha_core/n344_152 ),
	.I1(\top/processor/sha_core/n344_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_185 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s213  (
	.I0(\top/processor/sha_core/n344_154 ),
	.I1(\top/processor/sha_core/n344_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_187 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s214  (
	.I0(\top/processor/sha_core/n344_156 ),
	.I1(\top/processor/sha_core/n344_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_189 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s215  (
	.I0(\top/processor/sha_core/n344_158 ),
	.I1(\top/processor/sha_core/n344_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_191 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s216  (
	.I0(\top/processor/sha_core/n344_160 ),
	.I1(\top/processor/sha_core/n344_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_193 )
);
MUX2_LUT5 \top/processor/sha_core/n344_s217  (
	.I0(\top/processor/sha_core/n344_162 ),
	.I1(\top/processor/sha_core/n344_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n344_195 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s202  (
	.I0(\top/processor/sha_core/n345_132 ),
	.I1(\top/processor/sha_core/n345_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_165 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s203  (
	.I0(\top/processor/sha_core/n345_134 ),
	.I1(\top/processor/sha_core/n345_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_167 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s204  (
	.I0(\top/processor/sha_core/n345_136 ),
	.I1(\top/processor/sha_core/n345_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_169 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s205  (
	.I0(\top/processor/sha_core/n345_138 ),
	.I1(\top/processor/sha_core/n345_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_171 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s206  (
	.I0(\top/processor/sha_core/n345_140 ),
	.I1(\top/processor/sha_core/n345_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_173 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s207  (
	.I0(\top/processor/sha_core/n345_142 ),
	.I1(\top/processor/sha_core/n345_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_175 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s208  (
	.I0(\top/processor/sha_core/n345_144 ),
	.I1(\top/processor/sha_core/n345_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_177 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s209  (
	.I0(\top/processor/sha_core/n345_146 ),
	.I1(\top/processor/sha_core/n345_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_179 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s210  (
	.I0(\top/processor/sha_core/n345_148 ),
	.I1(\top/processor/sha_core/n345_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_181 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s211  (
	.I0(\top/processor/sha_core/n345_150 ),
	.I1(\top/processor/sha_core/n345_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_183 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s212  (
	.I0(\top/processor/sha_core/n345_152 ),
	.I1(\top/processor/sha_core/n345_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_185 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s213  (
	.I0(\top/processor/sha_core/n345_154 ),
	.I1(\top/processor/sha_core/n345_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_187 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s214  (
	.I0(\top/processor/sha_core/n345_156 ),
	.I1(\top/processor/sha_core/n345_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_189 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s215  (
	.I0(\top/processor/sha_core/n345_158 ),
	.I1(\top/processor/sha_core/n345_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_191 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s216  (
	.I0(\top/processor/sha_core/n345_160 ),
	.I1(\top/processor/sha_core/n345_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_193 )
);
MUX2_LUT5 \top/processor/sha_core/n345_s217  (
	.I0(\top/processor/sha_core/n345_162 ),
	.I1(\top/processor/sha_core/n345_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n345_195 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s202  (
	.I0(\top/processor/sha_core/n346_132 ),
	.I1(\top/processor/sha_core/n346_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_165 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s203  (
	.I0(\top/processor/sha_core/n346_134 ),
	.I1(\top/processor/sha_core/n346_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_167 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s204  (
	.I0(\top/processor/sha_core/n346_136 ),
	.I1(\top/processor/sha_core/n346_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_169 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s205  (
	.I0(\top/processor/sha_core/n346_138 ),
	.I1(\top/processor/sha_core/n346_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_171 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s206  (
	.I0(\top/processor/sha_core/n346_140 ),
	.I1(\top/processor/sha_core/n346_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_173 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s207  (
	.I0(\top/processor/sha_core/n346_142 ),
	.I1(\top/processor/sha_core/n346_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_175 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s208  (
	.I0(\top/processor/sha_core/n346_144 ),
	.I1(\top/processor/sha_core/n346_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_177 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s209  (
	.I0(\top/processor/sha_core/n346_146 ),
	.I1(\top/processor/sha_core/n346_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_179 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s210  (
	.I0(\top/processor/sha_core/n346_148 ),
	.I1(\top/processor/sha_core/n346_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_181 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s211  (
	.I0(\top/processor/sha_core/n346_150 ),
	.I1(\top/processor/sha_core/n346_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_183 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s212  (
	.I0(\top/processor/sha_core/n346_152 ),
	.I1(\top/processor/sha_core/n346_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_185 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s213  (
	.I0(\top/processor/sha_core/n346_154 ),
	.I1(\top/processor/sha_core/n346_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_187 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s214  (
	.I0(\top/processor/sha_core/n346_156 ),
	.I1(\top/processor/sha_core/n346_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_189 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s215  (
	.I0(\top/processor/sha_core/n346_158 ),
	.I1(\top/processor/sha_core/n346_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_191 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s216  (
	.I0(\top/processor/sha_core/n346_160 ),
	.I1(\top/processor/sha_core/n346_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_193 )
);
MUX2_LUT5 \top/processor/sha_core/n346_s217  (
	.I0(\top/processor/sha_core/n346_162 ),
	.I1(\top/processor/sha_core/n346_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n346_195 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s202  (
	.I0(\top/processor/sha_core/n347_132 ),
	.I1(\top/processor/sha_core/n347_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_165 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s203  (
	.I0(\top/processor/sha_core/n347_134 ),
	.I1(\top/processor/sha_core/n347_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_167 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s204  (
	.I0(\top/processor/sha_core/n347_136 ),
	.I1(\top/processor/sha_core/n347_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_169 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s205  (
	.I0(\top/processor/sha_core/n347_138 ),
	.I1(\top/processor/sha_core/n347_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_171 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s206  (
	.I0(\top/processor/sha_core/n347_140 ),
	.I1(\top/processor/sha_core/n347_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_173 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s207  (
	.I0(\top/processor/sha_core/n347_142 ),
	.I1(\top/processor/sha_core/n347_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_175 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s208  (
	.I0(\top/processor/sha_core/n347_144 ),
	.I1(\top/processor/sha_core/n347_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_177 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s209  (
	.I0(\top/processor/sha_core/n347_146 ),
	.I1(\top/processor/sha_core/n347_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_179 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s210  (
	.I0(\top/processor/sha_core/n347_148 ),
	.I1(\top/processor/sha_core/n347_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_181 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s211  (
	.I0(\top/processor/sha_core/n347_150 ),
	.I1(\top/processor/sha_core/n347_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_183 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s212  (
	.I0(\top/processor/sha_core/n347_152 ),
	.I1(\top/processor/sha_core/n347_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_185 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s213  (
	.I0(\top/processor/sha_core/n347_154 ),
	.I1(\top/processor/sha_core/n347_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_187 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s214  (
	.I0(\top/processor/sha_core/n347_156 ),
	.I1(\top/processor/sha_core/n347_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_189 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s215  (
	.I0(\top/processor/sha_core/n347_158 ),
	.I1(\top/processor/sha_core/n347_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_191 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s216  (
	.I0(\top/processor/sha_core/n347_160 ),
	.I1(\top/processor/sha_core/n347_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_193 )
);
MUX2_LUT5 \top/processor/sha_core/n347_s217  (
	.I0(\top/processor/sha_core/n347_162 ),
	.I1(\top/processor/sha_core/n347_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n347_195 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s202  (
	.I0(\top/processor/sha_core/n348_132 ),
	.I1(\top/processor/sha_core/n348_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_165 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s203  (
	.I0(\top/processor/sha_core/n348_134 ),
	.I1(\top/processor/sha_core/n348_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_167 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s204  (
	.I0(\top/processor/sha_core/n348_136 ),
	.I1(\top/processor/sha_core/n348_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_169 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s205  (
	.I0(\top/processor/sha_core/n348_138 ),
	.I1(\top/processor/sha_core/n348_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_171 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s206  (
	.I0(\top/processor/sha_core/n348_140 ),
	.I1(\top/processor/sha_core/n348_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_173 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s207  (
	.I0(\top/processor/sha_core/n348_142 ),
	.I1(\top/processor/sha_core/n348_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_175 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s208  (
	.I0(\top/processor/sha_core/n348_144 ),
	.I1(\top/processor/sha_core/n348_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_177 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s209  (
	.I0(\top/processor/sha_core/n348_146 ),
	.I1(\top/processor/sha_core/n348_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_179 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s210  (
	.I0(\top/processor/sha_core/n348_148 ),
	.I1(\top/processor/sha_core/n348_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_181 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s211  (
	.I0(\top/processor/sha_core/n348_150 ),
	.I1(\top/processor/sha_core/n348_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_183 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s212  (
	.I0(\top/processor/sha_core/n348_152 ),
	.I1(\top/processor/sha_core/n348_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_185 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s213  (
	.I0(\top/processor/sha_core/n348_154 ),
	.I1(\top/processor/sha_core/n348_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_187 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s214  (
	.I0(\top/processor/sha_core/n348_156 ),
	.I1(\top/processor/sha_core/n348_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_189 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s215  (
	.I0(\top/processor/sha_core/n348_158 ),
	.I1(\top/processor/sha_core/n348_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_191 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s216  (
	.I0(\top/processor/sha_core/n348_160 ),
	.I1(\top/processor/sha_core/n348_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_193 )
);
MUX2_LUT5 \top/processor/sha_core/n348_s217  (
	.I0(\top/processor/sha_core/n348_162 ),
	.I1(\top/processor/sha_core/n348_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n348_195 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s202  (
	.I0(\top/processor/sha_core/n349_132 ),
	.I1(\top/processor/sha_core/n349_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_165 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s203  (
	.I0(\top/processor/sha_core/n349_134 ),
	.I1(\top/processor/sha_core/n349_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_167 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s204  (
	.I0(\top/processor/sha_core/n349_136 ),
	.I1(\top/processor/sha_core/n349_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_169 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s205  (
	.I0(\top/processor/sha_core/n349_138 ),
	.I1(\top/processor/sha_core/n349_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_171 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s206  (
	.I0(\top/processor/sha_core/n349_140 ),
	.I1(\top/processor/sha_core/n349_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_173 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s207  (
	.I0(\top/processor/sha_core/n349_142 ),
	.I1(\top/processor/sha_core/n349_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_175 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s208  (
	.I0(\top/processor/sha_core/n349_144 ),
	.I1(\top/processor/sha_core/n349_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_177 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s209  (
	.I0(\top/processor/sha_core/n349_146 ),
	.I1(\top/processor/sha_core/n349_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_179 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s210  (
	.I0(\top/processor/sha_core/n349_148 ),
	.I1(\top/processor/sha_core/n349_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_181 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s211  (
	.I0(\top/processor/sha_core/n349_150 ),
	.I1(\top/processor/sha_core/n349_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_183 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s212  (
	.I0(\top/processor/sha_core/n349_152 ),
	.I1(\top/processor/sha_core/n349_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_185 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s213  (
	.I0(\top/processor/sha_core/n349_154 ),
	.I1(\top/processor/sha_core/n349_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_187 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s214  (
	.I0(\top/processor/sha_core/n349_156 ),
	.I1(\top/processor/sha_core/n349_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_189 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s215  (
	.I0(\top/processor/sha_core/n349_158 ),
	.I1(\top/processor/sha_core/n349_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_191 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s216  (
	.I0(\top/processor/sha_core/n349_160 ),
	.I1(\top/processor/sha_core/n349_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_193 )
);
MUX2_LUT5 \top/processor/sha_core/n349_s217  (
	.I0(\top/processor/sha_core/n349_162 ),
	.I1(\top/processor/sha_core/n349_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n349_195 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s202  (
	.I0(\top/processor/sha_core/n350_132 ),
	.I1(\top/processor/sha_core/n350_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_165 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s203  (
	.I0(\top/processor/sha_core/n350_134 ),
	.I1(\top/processor/sha_core/n350_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_167 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s204  (
	.I0(\top/processor/sha_core/n350_136 ),
	.I1(\top/processor/sha_core/n350_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_169 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s205  (
	.I0(\top/processor/sha_core/n350_138 ),
	.I1(\top/processor/sha_core/n350_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_171 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s206  (
	.I0(\top/processor/sha_core/n350_140 ),
	.I1(\top/processor/sha_core/n350_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_173 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s207  (
	.I0(\top/processor/sha_core/n350_142 ),
	.I1(\top/processor/sha_core/n350_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_175 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s208  (
	.I0(\top/processor/sha_core/n350_144 ),
	.I1(\top/processor/sha_core/n350_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_177 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s209  (
	.I0(\top/processor/sha_core/n350_146 ),
	.I1(\top/processor/sha_core/n350_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_179 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s210  (
	.I0(\top/processor/sha_core/n350_148 ),
	.I1(\top/processor/sha_core/n350_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_181 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s211  (
	.I0(\top/processor/sha_core/n350_150 ),
	.I1(\top/processor/sha_core/n350_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_183 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s212  (
	.I0(\top/processor/sha_core/n350_152 ),
	.I1(\top/processor/sha_core/n350_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_185 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s213  (
	.I0(\top/processor/sha_core/n350_154 ),
	.I1(\top/processor/sha_core/n350_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_187 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s214  (
	.I0(\top/processor/sha_core/n350_156 ),
	.I1(\top/processor/sha_core/n350_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_189 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s215  (
	.I0(\top/processor/sha_core/n350_158 ),
	.I1(\top/processor/sha_core/n350_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_191 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s216  (
	.I0(\top/processor/sha_core/n350_160 ),
	.I1(\top/processor/sha_core/n350_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_193 )
);
MUX2_LUT5 \top/processor/sha_core/n350_s217  (
	.I0(\top/processor/sha_core/n350_162 ),
	.I1(\top/processor/sha_core/n350_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n350_195 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s202  (
	.I0(\top/processor/sha_core/n351_132 ),
	.I1(\top/processor/sha_core/n351_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_165 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s203  (
	.I0(\top/processor/sha_core/n351_134 ),
	.I1(\top/processor/sha_core/n351_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_167 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s204  (
	.I0(\top/processor/sha_core/n351_136 ),
	.I1(\top/processor/sha_core/n351_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_169 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s205  (
	.I0(\top/processor/sha_core/n351_138 ),
	.I1(\top/processor/sha_core/n351_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_171 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s206  (
	.I0(\top/processor/sha_core/n351_140 ),
	.I1(\top/processor/sha_core/n351_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_173 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s207  (
	.I0(\top/processor/sha_core/n351_142 ),
	.I1(\top/processor/sha_core/n351_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_175 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s208  (
	.I0(\top/processor/sha_core/n351_144 ),
	.I1(\top/processor/sha_core/n351_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_177 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s209  (
	.I0(\top/processor/sha_core/n351_146 ),
	.I1(\top/processor/sha_core/n351_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_179 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s210  (
	.I0(\top/processor/sha_core/n351_148 ),
	.I1(\top/processor/sha_core/n351_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_181 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s211  (
	.I0(\top/processor/sha_core/n351_150 ),
	.I1(\top/processor/sha_core/n351_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_183 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s212  (
	.I0(\top/processor/sha_core/n351_152 ),
	.I1(\top/processor/sha_core/n351_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_185 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s213  (
	.I0(\top/processor/sha_core/n351_154 ),
	.I1(\top/processor/sha_core/n351_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_187 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s214  (
	.I0(\top/processor/sha_core/n351_156 ),
	.I1(\top/processor/sha_core/n351_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_189 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s215  (
	.I0(\top/processor/sha_core/n351_158 ),
	.I1(\top/processor/sha_core/n351_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_191 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s216  (
	.I0(\top/processor/sha_core/n351_160 ),
	.I1(\top/processor/sha_core/n351_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_193 )
);
MUX2_LUT5 \top/processor/sha_core/n351_s217  (
	.I0(\top/processor/sha_core/n351_162 ),
	.I1(\top/processor/sha_core/n351_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n351_195 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s202  (
	.I0(\top/processor/sha_core/n352_132 ),
	.I1(\top/processor/sha_core/n352_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_165 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s203  (
	.I0(\top/processor/sha_core/n352_134 ),
	.I1(\top/processor/sha_core/n352_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_167 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s204  (
	.I0(\top/processor/sha_core/n352_136 ),
	.I1(\top/processor/sha_core/n352_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_169 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s205  (
	.I0(\top/processor/sha_core/n352_138 ),
	.I1(\top/processor/sha_core/n352_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_171 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s206  (
	.I0(\top/processor/sha_core/n352_140 ),
	.I1(\top/processor/sha_core/n352_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_173 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s207  (
	.I0(\top/processor/sha_core/n352_142 ),
	.I1(\top/processor/sha_core/n352_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_175 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s208  (
	.I0(\top/processor/sha_core/n352_144 ),
	.I1(\top/processor/sha_core/n352_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_177 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s209  (
	.I0(\top/processor/sha_core/n352_146 ),
	.I1(\top/processor/sha_core/n352_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_179 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s210  (
	.I0(\top/processor/sha_core/n352_148 ),
	.I1(\top/processor/sha_core/n352_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_181 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s211  (
	.I0(\top/processor/sha_core/n352_150 ),
	.I1(\top/processor/sha_core/n352_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_183 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s212  (
	.I0(\top/processor/sha_core/n352_152 ),
	.I1(\top/processor/sha_core/n352_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_185 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s213  (
	.I0(\top/processor/sha_core/n352_154 ),
	.I1(\top/processor/sha_core/n352_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_187 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s214  (
	.I0(\top/processor/sha_core/n352_156 ),
	.I1(\top/processor/sha_core/n352_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_189 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s215  (
	.I0(\top/processor/sha_core/n352_158 ),
	.I1(\top/processor/sha_core/n352_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_191 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s216  (
	.I0(\top/processor/sha_core/n352_160 ),
	.I1(\top/processor/sha_core/n352_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_193 )
);
MUX2_LUT5 \top/processor/sha_core/n352_s217  (
	.I0(\top/processor/sha_core/n352_162 ),
	.I1(\top/processor/sha_core/n352_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n352_195 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s202  (
	.I0(\top/processor/sha_core/n353_132 ),
	.I1(\top/processor/sha_core/n353_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_165 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s203  (
	.I0(\top/processor/sha_core/n353_134 ),
	.I1(\top/processor/sha_core/n353_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_167 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s204  (
	.I0(\top/processor/sha_core/n353_136 ),
	.I1(\top/processor/sha_core/n353_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_169 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s205  (
	.I0(\top/processor/sha_core/n353_138 ),
	.I1(\top/processor/sha_core/n353_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_171 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s206  (
	.I0(\top/processor/sha_core/n353_140 ),
	.I1(\top/processor/sha_core/n353_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_173 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s207  (
	.I0(\top/processor/sha_core/n353_142 ),
	.I1(\top/processor/sha_core/n353_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_175 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s208  (
	.I0(\top/processor/sha_core/n353_144 ),
	.I1(\top/processor/sha_core/n353_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_177 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s209  (
	.I0(\top/processor/sha_core/n353_146 ),
	.I1(\top/processor/sha_core/n353_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_179 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s210  (
	.I0(\top/processor/sha_core/n353_148 ),
	.I1(\top/processor/sha_core/n353_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_181 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s211  (
	.I0(\top/processor/sha_core/n353_150 ),
	.I1(\top/processor/sha_core/n353_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_183 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s212  (
	.I0(\top/processor/sha_core/n353_152 ),
	.I1(\top/processor/sha_core/n353_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_185 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s213  (
	.I0(\top/processor/sha_core/n353_154 ),
	.I1(\top/processor/sha_core/n353_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_187 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s214  (
	.I0(\top/processor/sha_core/n353_156 ),
	.I1(\top/processor/sha_core/n353_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_189 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s215  (
	.I0(\top/processor/sha_core/n353_158 ),
	.I1(\top/processor/sha_core/n353_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_191 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s216  (
	.I0(\top/processor/sha_core/n353_160 ),
	.I1(\top/processor/sha_core/n353_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_193 )
);
MUX2_LUT5 \top/processor/sha_core/n353_s217  (
	.I0(\top/processor/sha_core/n353_162 ),
	.I1(\top/processor/sha_core/n353_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n353_195 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s202  (
	.I0(\top/processor/sha_core/n354_132 ),
	.I1(\top/processor/sha_core/n354_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_165 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s203  (
	.I0(\top/processor/sha_core/n354_134 ),
	.I1(\top/processor/sha_core/n354_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_167 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s204  (
	.I0(\top/processor/sha_core/n354_136 ),
	.I1(\top/processor/sha_core/n354_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_169 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s205  (
	.I0(\top/processor/sha_core/n354_138 ),
	.I1(\top/processor/sha_core/n354_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_171 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s206  (
	.I0(\top/processor/sha_core/n354_140 ),
	.I1(\top/processor/sha_core/n354_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_173 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s207  (
	.I0(\top/processor/sha_core/n354_142 ),
	.I1(\top/processor/sha_core/n354_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_175 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s208  (
	.I0(\top/processor/sha_core/n354_144 ),
	.I1(\top/processor/sha_core/n354_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_177 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s209  (
	.I0(\top/processor/sha_core/n354_146 ),
	.I1(\top/processor/sha_core/n354_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_179 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s210  (
	.I0(\top/processor/sha_core/n354_148 ),
	.I1(\top/processor/sha_core/n354_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_181 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s211  (
	.I0(\top/processor/sha_core/n354_150 ),
	.I1(\top/processor/sha_core/n354_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_183 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s212  (
	.I0(\top/processor/sha_core/n354_152 ),
	.I1(\top/processor/sha_core/n354_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_185 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s213  (
	.I0(\top/processor/sha_core/n354_154 ),
	.I1(\top/processor/sha_core/n354_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_187 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s214  (
	.I0(\top/processor/sha_core/n354_156 ),
	.I1(\top/processor/sha_core/n354_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_189 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s215  (
	.I0(\top/processor/sha_core/n354_158 ),
	.I1(\top/processor/sha_core/n354_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_191 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s216  (
	.I0(\top/processor/sha_core/n354_160 ),
	.I1(\top/processor/sha_core/n354_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_193 )
);
MUX2_LUT5 \top/processor/sha_core/n354_s217  (
	.I0(\top/processor/sha_core/n354_162 ),
	.I1(\top/processor/sha_core/n354_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n354_195 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s202  (
	.I0(\top/processor/sha_core/n355_132 ),
	.I1(\top/processor/sha_core/n355_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_165 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s203  (
	.I0(\top/processor/sha_core/n355_134 ),
	.I1(\top/processor/sha_core/n355_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_167 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s204  (
	.I0(\top/processor/sha_core/n355_136 ),
	.I1(\top/processor/sha_core/n355_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_169 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s205  (
	.I0(\top/processor/sha_core/n355_138 ),
	.I1(\top/processor/sha_core/n355_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_171 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s206  (
	.I0(\top/processor/sha_core/n355_140 ),
	.I1(\top/processor/sha_core/n355_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_173 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s207  (
	.I0(\top/processor/sha_core/n355_142 ),
	.I1(\top/processor/sha_core/n355_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_175 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s208  (
	.I0(\top/processor/sha_core/n355_144 ),
	.I1(\top/processor/sha_core/n355_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_177 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s209  (
	.I0(\top/processor/sha_core/n355_146 ),
	.I1(\top/processor/sha_core/n355_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_179 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s210  (
	.I0(\top/processor/sha_core/n355_148 ),
	.I1(\top/processor/sha_core/n355_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_181 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s211  (
	.I0(\top/processor/sha_core/n355_150 ),
	.I1(\top/processor/sha_core/n355_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_183 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s212  (
	.I0(\top/processor/sha_core/n355_152 ),
	.I1(\top/processor/sha_core/n355_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_185 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s213  (
	.I0(\top/processor/sha_core/n355_154 ),
	.I1(\top/processor/sha_core/n355_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_187 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s214  (
	.I0(\top/processor/sha_core/n355_156 ),
	.I1(\top/processor/sha_core/n355_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_189 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s215  (
	.I0(\top/processor/sha_core/n355_158 ),
	.I1(\top/processor/sha_core/n355_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_191 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s216  (
	.I0(\top/processor/sha_core/n355_160 ),
	.I1(\top/processor/sha_core/n355_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_193 )
);
MUX2_LUT5 \top/processor/sha_core/n355_s217  (
	.I0(\top/processor/sha_core/n355_162 ),
	.I1(\top/processor/sha_core/n355_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n355_195 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s202  (
	.I0(\top/processor/sha_core/n356_132 ),
	.I1(\top/processor/sha_core/n356_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_165 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s203  (
	.I0(\top/processor/sha_core/n356_134 ),
	.I1(\top/processor/sha_core/n356_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_167 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s204  (
	.I0(\top/processor/sha_core/n356_136 ),
	.I1(\top/processor/sha_core/n356_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_169 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s205  (
	.I0(\top/processor/sha_core/n356_138 ),
	.I1(\top/processor/sha_core/n356_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_171 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s206  (
	.I0(\top/processor/sha_core/n356_140 ),
	.I1(\top/processor/sha_core/n356_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_173 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s207  (
	.I0(\top/processor/sha_core/n356_142 ),
	.I1(\top/processor/sha_core/n356_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_175 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s208  (
	.I0(\top/processor/sha_core/n356_144 ),
	.I1(\top/processor/sha_core/n356_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_177 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s209  (
	.I0(\top/processor/sha_core/n356_146 ),
	.I1(\top/processor/sha_core/n356_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_179 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s210  (
	.I0(\top/processor/sha_core/n356_148 ),
	.I1(\top/processor/sha_core/n356_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_181 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s211  (
	.I0(\top/processor/sha_core/n356_150 ),
	.I1(\top/processor/sha_core/n356_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_183 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s212  (
	.I0(\top/processor/sha_core/n356_152 ),
	.I1(\top/processor/sha_core/n356_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_185 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s213  (
	.I0(\top/processor/sha_core/n356_154 ),
	.I1(\top/processor/sha_core/n356_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_187 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s214  (
	.I0(\top/processor/sha_core/n356_156 ),
	.I1(\top/processor/sha_core/n356_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_189 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s215  (
	.I0(\top/processor/sha_core/n356_158 ),
	.I1(\top/processor/sha_core/n356_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_191 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s216  (
	.I0(\top/processor/sha_core/n356_160 ),
	.I1(\top/processor/sha_core/n356_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_193 )
);
MUX2_LUT5 \top/processor/sha_core/n356_s217  (
	.I0(\top/processor/sha_core/n356_162 ),
	.I1(\top/processor/sha_core/n356_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n356_195 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s202  (
	.I0(\top/processor/sha_core/n357_132 ),
	.I1(\top/processor/sha_core/n357_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_165 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s203  (
	.I0(\top/processor/sha_core/n357_134 ),
	.I1(\top/processor/sha_core/n357_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_167 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s204  (
	.I0(\top/processor/sha_core/n357_136 ),
	.I1(\top/processor/sha_core/n357_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_169 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s205  (
	.I0(\top/processor/sha_core/n357_138 ),
	.I1(\top/processor/sha_core/n357_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_171 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s206  (
	.I0(\top/processor/sha_core/n357_140 ),
	.I1(\top/processor/sha_core/n357_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_173 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s207  (
	.I0(\top/processor/sha_core/n357_142 ),
	.I1(\top/processor/sha_core/n357_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_175 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s208  (
	.I0(\top/processor/sha_core/n357_144 ),
	.I1(\top/processor/sha_core/n357_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_177 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s209  (
	.I0(\top/processor/sha_core/n357_146 ),
	.I1(\top/processor/sha_core/n357_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_179 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s210  (
	.I0(\top/processor/sha_core/n357_148 ),
	.I1(\top/processor/sha_core/n357_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_181 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s211  (
	.I0(\top/processor/sha_core/n357_150 ),
	.I1(\top/processor/sha_core/n357_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_183 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s212  (
	.I0(\top/processor/sha_core/n357_152 ),
	.I1(\top/processor/sha_core/n357_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_185 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s213  (
	.I0(\top/processor/sha_core/n357_154 ),
	.I1(\top/processor/sha_core/n357_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_187 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s214  (
	.I0(\top/processor/sha_core/n357_156 ),
	.I1(\top/processor/sha_core/n357_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_189 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s215  (
	.I0(\top/processor/sha_core/n357_158 ),
	.I1(\top/processor/sha_core/n357_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_191 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s216  (
	.I0(\top/processor/sha_core/n357_160 ),
	.I1(\top/processor/sha_core/n357_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_193 )
);
MUX2_LUT5 \top/processor/sha_core/n357_s217  (
	.I0(\top/processor/sha_core/n357_162 ),
	.I1(\top/processor/sha_core/n357_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n357_195 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s202  (
	.I0(\top/processor/sha_core/n358_132 ),
	.I1(\top/processor/sha_core/n358_133 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_165 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s203  (
	.I0(\top/processor/sha_core/n358_134 ),
	.I1(\top/processor/sha_core/n358_135 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_167 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s204  (
	.I0(\top/processor/sha_core/n358_136 ),
	.I1(\top/processor/sha_core/n358_137 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_169 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s205  (
	.I0(\top/processor/sha_core/n358_138 ),
	.I1(\top/processor/sha_core/n358_139 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_171 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s206  (
	.I0(\top/processor/sha_core/n358_140 ),
	.I1(\top/processor/sha_core/n358_141 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_173 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s207  (
	.I0(\top/processor/sha_core/n358_142 ),
	.I1(\top/processor/sha_core/n358_143 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_175 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s208  (
	.I0(\top/processor/sha_core/n358_144 ),
	.I1(\top/processor/sha_core/n358_145 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_177 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s209  (
	.I0(\top/processor/sha_core/n358_146 ),
	.I1(\top/processor/sha_core/n358_147 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_179 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s210  (
	.I0(\top/processor/sha_core/n358_148 ),
	.I1(\top/processor/sha_core/n358_149 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_181 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s211  (
	.I0(\top/processor/sha_core/n358_150 ),
	.I1(\top/processor/sha_core/n358_151 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_183 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s212  (
	.I0(\top/processor/sha_core/n358_152 ),
	.I1(\top/processor/sha_core/n358_153 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_185 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s213  (
	.I0(\top/processor/sha_core/n358_154 ),
	.I1(\top/processor/sha_core/n358_155 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_187 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s214  (
	.I0(\top/processor/sha_core/n358_156 ),
	.I1(\top/processor/sha_core/n358_157 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_189 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s215  (
	.I0(\top/processor/sha_core/n358_158 ),
	.I1(\top/processor/sha_core/n358_159 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_191 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s216  (
	.I0(\top/processor/sha_core/n358_160 ),
	.I1(\top/processor/sha_core/n358_161 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_193 )
);
MUX2_LUT5 \top/processor/sha_core/n358_s217  (
	.I0(\top/processor/sha_core/n358_162 ),
	.I1(\top/processor/sha_core/n358_163 ),
	.S0(\top/processor/sha_core/t [1]),
	.O(\top/processor/sha_core/n358_195 )
);
MUX2_LUT5 \top/processor/sha_core/n3488_s176  (
	.I0(\top/processor/sha_core/n3488_139 ),
	.I1(\top/processor/sha_core/n3488_141 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3488_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3488_s177  (
	.I0(\top/processor/sha_core/n3488_143 ),
	.I1(\top/processor/sha_core/n3488_145 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3488_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3488_s178  (
	.I0(\top/processor/sha_core/n3488_147 ),
	.I1(\top/processor/sha_core/n3488_133 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3488_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3488_s179  (
	.I0(\top/processor/sha_core/n3488_135 ),
	.I1(\top/processor/sha_core/n3488_137 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3488_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3489_s176  (
	.I0(\top/processor/sha_core/n3489_133 ),
	.I1(\top/processor/sha_core/n3489_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3489_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3489_s177  (
	.I0(\top/processor/sha_core/n3489_137 ),
	.I1(\top/processor/sha_core/n3489_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3489_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3489_s178  (
	.I0(\top/processor/sha_core/n3489_141 ),
	.I1(\top/processor/sha_core/n3489_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3489_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3489_s179  (
	.I0(\top/processor/sha_core/n3489_145 ),
	.I1(\top/processor/sha_core/n3489_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3489_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3490_s176  (
	.I0(\top/processor/sha_core/n3490_133 ),
	.I1(\top/processor/sha_core/n3490_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3490_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3490_s177  (
	.I0(\top/processor/sha_core/n3490_137 ),
	.I1(\top/processor/sha_core/n3490_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3490_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3490_s178  (
	.I0(\top/processor/sha_core/n3490_141 ),
	.I1(\top/processor/sha_core/n3490_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3490_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3490_s179  (
	.I0(\top/processor/sha_core/n3490_145 ),
	.I1(\top/processor/sha_core/n3490_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3490_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3491_s176  (
	.I0(\top/processor/sha_core/n3491_133 ),
	.I1(\top/processor/sha_core/n3491_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3491_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3491_s177  (
	.I0(\top/processor/sha_core/n3491_137 ),
	.I1(\top/processor/sha_core/n3491_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3491_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3491_s178  (
	.I0(\top/processor/sha_core/n3491_141 ),
	.I1(\top/processor/sha_core/n3491_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3491_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3491_s179  (
	.I0(\top/processor/sha_core/n3491_145 ),
	.I1(\top/processor/sha_core/n3491_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3491_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3492_s176  (
	.I0(\top/processor/sha_core/n3492_133 ),
	.I1(\top/processor/sha_core/n3492_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3492_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3492_s177  (
	.I0(\top/processor/sha_core/n3492_137 ),
	.I1(\top/processor/sha_core/n3492_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3492_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3492_s178  (
	.I0(\top/processor/sha_core/n3492_141 ),
	.I1(\top/processor/sha_core/n3492_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3492_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3492_s179  (
	.I0(\top/processor/sha_core/n3492_145 ),
	.I1(\top/processor/sha_core/n3492_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3492_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3493_s176  (
	.I0(\top/processor/sha_core/n3493_133 ),
	.I1(\top/processor/sha_core/n3493_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3493_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3493_s177  (
	.I0(\top/processor/sha_core/n3493_137 ),
	.I1(\top/processor/sha_core/n3493_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3493_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3493_s178  (
	.I0(\top/processor/sha_core/n3493_141 ),
	.I1(\top/processor/sha_core/n3493_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3493_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3493_s179  (
	.I0(\top/processor/sha_core/n3493_145 ),
	.I1(\top/processor/sha_core/n3493_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3493_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3494_s176  (
	.I0(\top/processor/sha_core/n3494_145 ),
	.I1(\top/processor/sha_core/n3494_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3494_182 )
);
MUX2_LUT5 \top/processor/sha_core/n3494_s177  (
	.I0(\top/processor/sha_core/n3494_148 ),
	.I1(\top/processor/sha_core/n3494_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3494_184 )
);
MUX2_LUT5 \top/processor/sha_core/n3494_s178  (
	.I0(\top/processor/sha_core/n3494_137 ),
	.I1(\top/processor/sha_core/n3494_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3494_186 )
);
MUX2_LUT5 \top/processor/sha_core/n3494_s179  (
	.I0(\top/processor/sha_core/n3494_141 ),
	.I1(\top/processor/sha_core/n3494_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3494_188 )
);
MUX2_LUT5 \top/processor/sha_core/n3495_s176  (
	.I0(\top/processor/sha_core/n3495_133 ),
	.I1(\top/processor/sha_core/n3495_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3495_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3495_s177  (
	.I0(\top/processor/sha_core/n3495_137 ),
	.I1(\top/processor/sha_core/n3495_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3495_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3495_s178  (
	.I0(\top/processor/sha_core/n3495_141 ),
	.I1(\top/processor/sha_core/n3495_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3495_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3495_s179  (
	.I0(\top/processor/sha_core/n3495_145 ),
	.I1(\top/processor/sha_core/n3495_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3495_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3496_s176  (
	.I0(\top/processor/sha_core/n3496_133 ),
	.I1(\top/processor/sha_core/n3496_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3496_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3496_s177  (
	.I0(\top/processor/sha_core/n3496_137 ),
	.I1(\top/processor/sha_core/n3496_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3496_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3496_s178  (
	.I0(\top/processor/sha_core/n3496_141 ),
	.I1(\top/processor/sha_core/n3496_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3496_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3496_s179  (
	.I0(\top/processor/sha_core/n3496_145 ),
	.I1(\top/processor/sha_core/n3496_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3496_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3497_s176  (
	.I0(\top/processor/sha_core/n3497_133 ),
	.I1(\top/processor/sha_core/n3497_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3497_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3497_s177  (
	.I0(\top/processor/sha_core/n3497_137 ),
	.I1(\top/processor/sha_core/n3497_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3497_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3497_s178  (
	.I0(\top/processor/sha_core/n3497_141 ),
	.I1(\top/processor/sha_core/n3497_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3497_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3497_s179  (
	.I0(\top/processor/sha_core/n3497_145 ),
	.I1(\top/processor/sha_core/n3497_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3497_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3498_s176  (
	.I0(\top/processor/sha_core/n3498_133 ),
	.I1(\top/processor/sha_core/n3498_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3498_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3498_s177  (
	.I0(\top/processor/sha_core/n3498_137 ),
	.I1(\top/processor/sha_core/n3498_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3498_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3498_s178  (
	.I0(\top/processor/sha_core/n3498_141 ),
	.I1(\top/processor/sha_core/n3498_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3498_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3498_s179  (
	.I0(\top/processor/sha_core/n3498_145 ),
	.I1(\top/processor/sha_core/n3498_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3498_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3499_s176  (
	.I0(\top/processor/sha_core/n3499_133 ),
	.I1(\top/processor/sha_core/n3499_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3499_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3499_s177  (
	.I0(\top/processor/sha_core/n3499_137 ),
	.I1(\top/processor/sha_core/n3499_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3499_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3499_s178  (
	.I0(\top/processor/sha_core/n3499_141 ),
	.I1(\top/processor/sha_core/n3499_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3499_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3499_s179  (
	.I0(\top/processor/sha_core/n3499_145 ),
	.I1(\top/processor/sha_core/n3499_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3499_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3500_s176  (
	.I0(\top/processor/sha_core/n3500_133 ),
	.I1(\top/processor/sha_core/n3500_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3500_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3500_s177  (
	.I0(\top/processor/sha_core/n3500_137 ),
	.I1(\top/processor/sha_core/n3500_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3500_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3500_s178  (
	.I0(\top/processor/sha_core/n3500_141 ),
	.I1(\top/processor/sha_core/n3500_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3500_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3500_s179  (
	.I0(\top/processor/sha_core/n3500_145 ),
	.I1(\top/processor/sha_core/n3500_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3500_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3501_s176  (
	.I0(\top/processor/sha_core/n3501_133 ),
	.I1(\top/processor/sha_core/n3501_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3501_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3501_s177  (
	.I0(\top/processor/sha_core/n3501_137 ),
	.I1(\top/processor/sha_core/n3501_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3501_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3501_s178  (
	.I0(\top/processor/sha_core/n3501_141 ),
	.I1(\top/processor/sha_core/n3501_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3501_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3501_s179  (
	.I0(\top/processor/sha_core/n3501_145 ),
	.I1(\top/processor/sha_core/n3501_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3501_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3502_s176  (
	.I0(\top/processor/sha_core/n3502_133 ),
	.I1(\top/processor/sha_core/n3502_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3502_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3502_s177  (
	.I0(\top/processor/sha_core/n3502_137 ),
	.I1(\top/processor/sha_core/n3502_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3502_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3502_s178  (
	.I0(\top/processor/sha_core/n3502_141 ),
	.I1(\top/processor/sha_core/n3502_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3502_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3502_s179  (
	.I0(\top/processor/sha_core/n3502_145 ),
	.I1(\top/processor/sha_core/n3502_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3502_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3503_s176  (
	.I0(\top/processor/sha_core/n3503_133 ),
	.I1(\top/processor/sha_core/n3503_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3503_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3503_s177  (
	.I0(\top/processor/sha_core/n3503_137 ),
	.I1(\top/processor/sha_core/n3503_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3503_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3503_s178  (
	.I0(\top/processor/sha_core/n3503_141 ),
	.I1(\top/processor/sha_core/n3503_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3503_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3503_s179  (
	.I0(\top/processor/sha_core/n3503_145 ),
	.I1(\top/processor/sha_core/n3503_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3503_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3504_s176  (
	.I0(\top/processor/sha_core/n3504_133 ),
	.I1(\top/processor/sha_core/n3504_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3504_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3504_s177  (
	.I0(\top/processor/sha_core/n3504_137 ),
	.I1(\top/processor/sha_core/n3504_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3504_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3504_s178  (
	.I0(\top/processor/sha_core/n3504_141 ),
	.I1(\top/processor/sha_core/n3504_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3504_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3504_s179  (
	.I0(\top/processor/sha_core/n3504_145 ),
	.I1(\top/processor/sha_core/n3504_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3504_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3505_s176  (
	.I0(\top/processor/sha_core/n3505_133 ),
	.I1(\top/processor/sha_core/n3505_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3505_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3505_s177  (
	.I0(\top/processor/sha_core/n3505_137 ),
	.I1(\top/processor/sha_core/n3505_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3505_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3505_s178  (
	.I0(\top/processor/sha_core/n3505_141 ),
	.I1(\top/processor/sha_core/n3505_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3505_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3505_s179  (
	.I0(\top/processor/sha_core/n3505_145 ),
	.I1(\top/processor/sha_core/n3505_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3505_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3506_s176  (
	.I0(\top/processor/sha_core/n3506_133 ),
	.I1(\top/processor/sha_core/n3506_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3506_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3506_s177  (
	.I0(\top/processor/sha_core/n3506_137 ),
	.I1(\top/processor/sha_core/n3506_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3506_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3506_s178  (
	.I0(\top/processor/sha_core/n3506_141 ),
	.I1(\top/processor/sha_core/n3506_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3506_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3506_s179  (
	.I0(\top/processor/sha_core/n3506_145 ),
	.I1(\top/processor/sha_core/n3506_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3506_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3507_s176  (
	.I0(\top/processor/sha_core/n3507_133 ),
	.I1(\top/processor/sha_core/n3507_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3507_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3507_s177  (
	.I0(\top/processor/sha_core/n3507_137 ),
	.I1(\top/processor/sha_core/n3507_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3507_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3507_s178  (
	.I0(\top/processor/sha_core/n3507_141 ),
	.I1(\top/processor/sha_core/n3507_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3507_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3507_s179  (
	.I0(\top/processor/sha_core/n3507_145 ),
	.I1(\top/processor/sha_core/n3507_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3507_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3508_s176  (
	.I0(\top/processor/sha_core/n3508_133 ),
	.I1(\top/processor/sha_core/n3508_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3508_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3508_s177  (
	.I0(\top/processor/sha_core/n3508_137 ),
	.I1(\top/processor/sha_core/n3508_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3508_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3508_s178  (
	.I0(\top/processor/sha_core/n3508_141 ),
	.I1(\top/processor/sha_core/n3508_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3508_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3508_s179  (
	.I0(\top/processor/sha_core/n3508_145 ),
	.I1(\top/processor/sha_core/n3508_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3508_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3509_s176  (
	.I0(\top/processor/sha_core/n3509_133 ),
	.I1(\top/processor/sha_core/n3509_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3509_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3509_s177  (
	.I0(\top/processor/sha_core/n3509_137 ),
	.I1(\top/processor/sha_core/n3509_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3509_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3509_s178  (
	.I0(\top/processor/sha_core/n3509_141 ),
	.I1(\top/processor/sha_core/n3509_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3509_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3509_s179  (
	.I0(\top/processor/sha_core/n3509_145 ),
	.I1(\top/processor/sha_core/n3509_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3509_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3510_s176  (
	.I0(\top/processor/sha_core/n3510_133 ),
	.I1(\top/processor/sha_core/n3510_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3510_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3510_s177  (
	.I0(\top/processor/sha_core/n3510_137 ),
	.I1(\top/processor/sha_core/n3510_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3510_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3510_s178  (
	.I0(\top/processor/sha_core/n3510_141 ),
	.I1(\top/processor/sha_core/n3510_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3510_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3510_s179  (
	.I0(\top/processor/sha_core/n3510_145 ),
	.I1(\top/processor/sha_core/n3510_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3510_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3511_s176  (
	.I0(\top/processor/sha_core/n3511_133 ),
	.I1(\top/processor/sha_core/n3511_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3511_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3511_s177  (
	.I0(\top/processor/sha_core/n3511_137 ),
	.I1(\top/processor/sha_core/n3511_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3511_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3511_s178  (
	.I0(\top/processor/sha_core/n3511_141 ),
	.I1(\top/processor/sha_core/n3511_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3511_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3511_s179  (
	.I0(\top/processor/sha_core/n3511_145 ),
	.I1(\top/processor/sha_core/n3511_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3511_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3512_s176  (
	.I0(\top/processor/sha_core/n3512_133 ),
	.I1(\top/processor/sha_core/n3512_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3512_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3512_s177  (
	.I0(\top/processor/sha_core/n3512_137 ),
	.I1(\top/processor/sha_core/n3512_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3512_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3512_s178  (
	.I0(\top/processor/sha_core/n3512_141 ),
	.I1(\top/processor/sha_core/n3512_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3512_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3512_s179  (
	.I0(\top/processor/sha_core/n3512_145 ),
	.I1(\top/processor/sha_core/n3512_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3512_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3513_s176  (
	.I0(\top/processor/sha_core/n3513_133 ),
	.I1(\top/processor/sha_core/n3513_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3513_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3513_s177  (
	.I0(\top/processor/sha_core/n3513_137 ),
	.I1(\top/processor/sha_core/n3513_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3513_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3513_s178  (
	.I0(\top/processor/sha_core/n3513_141 ),
	.I1(\top/processor/sha_core/n3513_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3513_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3513_s179  (
	.I0(\top/processor/sha_core/n3513_145 ),
	.I1(\top/processor/sha_core/n3513_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3513_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3514_s176  (
	.I0(\top/processor/sha_core/n3514_133 ),
	.I1(\top/processor/sha_core/n3514_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3514_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3514_s177  (
	.I0(\top/processor/sha_core/n3514_137 ),
	.I1(\top/processor/sha_core/n3514_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3514_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3514_s178  (
	.I0(\top/processor/sha_core/n3514_141 ),
	.I1(\top/processor/sha_core/n3514_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3514_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3514_s179  (
	.I0(\top/processor/sha_core/n3514_145 ),
	.I1(\top/processor/sha_core/n3514_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3514_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3515_s176  (
	.I0(\top/processor/sha_core/n3515_133 ),
	.I1(\top/processor/sha_core/n3515_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3515_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3515_s177  (
	.I0(\top/processor/sha_core/n3515_137 ),
	.I1(\top/processor/sha_core/n3515_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3515_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3515_s178  (
	.I0(\top/processor/sha_core/n3515_141 ),
	.I1(\top/processor/sha_core/n3515_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3515_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3515_s179  (
	.I0(\top/processor/sha_core/n3515_145 ),
	.I1(\top/processor/sha_core/n3515_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3515_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3516_s176  (
	.I0(\top/processor/sha_core/n3516_133 ),
	.I1(\top/processor/sha_core/n3516_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3516_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3516_s177  (
	.I0(\top/processor/sha_core/n3516_137 ),
	.I1(\top/processor/sha_core/n3516_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3516_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3516_s178  (
	.I0(\top/processor/sha_core/n3516_141 ),
	.I1(\top/processor/sha_core/n3516_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3516_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3516_s179  (
	.I0(\top/processor/sha_core/n3516_145 ),
	.I1(\top/processor/sha_core/n3516_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3516_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3517_s176  (
	.I0(\top/processor/sha_core/n3517_133 ),
	.I1(\top/processor/sha_core/n3517_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3517_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3517_s177  (
	.I0(\top/processor/sha_core/n3517_137 ),
	.I1(\top/processor/sha_core/n3517_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3517_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3517_s178  (
	.I0(\top/processor/sha_core/n3517_141 ),
	.I1(\top/processor/sha_core/n3517_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3517_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3517_s179  (
	.I0(\top/processor/sha_core/n3517_145 ),
	.I1(\top/processor/sha_core/n3517_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3517_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3518_s176  (
	.I0(\top/processor/sha_core/n3518_133 ),
	.I1(\top/processor/sha_core/n3518_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3518_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3518_s177  (
	.I0(\top/processor/sha_core/n3518_137 ),
	.I1(\top/processor/sha_core/n3518_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3518_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3518_s178  (
	.I0(\top/processor/sha_core/n3518_141 ),
	.I1(\top/processor/sha_core/n3518_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3518_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3518_s179  (
	.I0(\top/processor/sha_core/n3518_145 ),
	.I1(\top/processor/sha_core/n3518_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3518_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3519_s176  (
	.I0(\top/processor/sha_core/n3519_133 ),
	.I1(\top/processor/sha_core/n3519_135 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3519_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3519_s177  (
	.I0(\top/processor/sha_core/n3519_137 ),
	.I1(\top/processor/sha_core/n3519_139 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3519_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3519_s178  (
	.I0(\top/processor/sha_core/n3519_141 ),
	.I1(\top/processor/sha_core/n3519_143 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3519_185 )
);
MUX2_LUT5 \top/processor/sha_core/n3519_s179  (
	.I0(\top/processor/sha_core/n3519_145 ),
	.I1(\top/processor/sha_core/n3519_147 ),
	.S0(\top/processor/sha_core/n3461_11 ),
	.O(\top/processor/sha_core/n3519_187 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s127  (
	.I0(\top/processor/sha_core/n3607_149 ),
	.I1(\top/processor/sha_core/n3607_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s128  (
	.I0(\top/processor/sha_core/n3607_153 ),
	.I1(\top/processor/sha_core/n3607_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s129  (
	.I0(\top/processor/sha_core/n3607_157 ),
	.I1(\top/processor/sha_core/n3607_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s130  (
	.I0(\top/processor/sha_core/n3607_161 ),
	.I1(\top/processor/sha_core/n3607_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s131  (
	.I0(\top/processor/sha_core/n3607_133 ),
	.I1(\top/processor/sha_core/n3607_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s132  (
	.I0(\top/processor/sha_core/n3607_137 ),
	.I1(\top/processor/sha_core/n3607_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s133  (
	.I0(\top/processor/sha_core/n3607_141 ),
	.I1(\top/processor/sha_core/n3607_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3705_s134  (
	.I0(\top/processor/sha_core/n3607_145 ),
	.I1(\top/processor/sha_core/n3607_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3705_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s127  (
	.I0(\top/processor/sha_core/n3608_149 ),
	.I1(\top/processor/sha_core/n3608_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s128  (
	.I0(\top/processor/sha_core/n3608_153 ),
	.I1(\top/processor/sha_core/n3608_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s129  (
	.I0(\top/processor/sha_core/n3608_157 ),
	.I1(\top/processor/sha_core/n3608_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s130  (
	.I0(\top/processor/sha_core/n3608_161 ),
	.I1(\top/processor/sha_core/n3608_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s131  (
	.I0(\top/processor/sha_core/n3608_133 ),
	.I1(\top/processor/sha_core/n3608_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s132  (
	.I0(\top/processor/sha_core/n3608_137 ),
	.I1(\top/processor/sha_core/n3608_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s133  (
	.I0(\top/processor/sha_core/n3608_141 ),
	.I1(\top/processor/sha_core/n3608_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3706_s134  (
	.I0(\top/processor/sha_core/n3608_145 ),
	.I1(\top/processor/sha_core/n3608_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3706_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s127  (
	.I0(\top/processor/sha_core/n3609_149 ),
	.I1(\top/processor/sha_core/n3609_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s128  (
	.I0(\top/processor/sha_core/n3609_153 ),
	.I1(\top/processor/sha_core/n3609_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s129  (
	.I0(\top/processor/sha_core/n3609_157 ),
	.I1(\top/processor/sha_core/n3609_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s130  (
	.I0(\top/processor/sha_core/n3609_161 ),
	.I1(\top/processor/sha_core/n3609_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s131  (
	.I0(\top/processor/sha_core/n3609_133 ),
	.I1(\top/processor/sha_core/n3609_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s132  (
	.I0(\top/processor/sha_core/n3609_137 ),
	.I1(\top/processor/sha_core/n3609_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s133  (
	.I0(\top/processor/sha_core/n3609_141 ),
	.I1(\top/processor/sha_core/n3609_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3707_s134  (
	.I0(\top/processor/sha_core/n3609_145 ),
	.I1(\top/processor/sha_core/n3609_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3707_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s127  (
	.I0(\top/processor/sha_core/n3610_149 ),
	.I1(\top/processor/sha_core/n3610_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s128  (
	.I0(\top/processor/sha_core/n3610_153 ),
	.I1(\top/processor/sha_core/n3610_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s129  (
	.I0(\top/processor/sha_core/n3610_157 ),
	.I1(\top/processor/sha_core/n3610_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s130  (
	.I0(\top/processor/sha_core/n3610_161 ),
	.I1(\top/processor/sha_core/n3610_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s131  (
	.I0(\top/processor/sha_core/n3610_133 ),
	.I1(\top/processor/sha_core/n3610_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s132  (
	.I0(\top/processor/sha_core/n3610_137 ),
	.I1(\top/processor/sha_core/n3610_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s133  (
	.I0(\top/processor/sha_core/n3610_141 ),
	.I1(\top/processor/sha_core/n3610_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3708_s134  (
	.I0(\top/processor/sha_core/n3610_145 ),
	.I1(\top/processor/sha_core/n3610_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3708_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s127  (
	.I0(\top/processor/sha_core/n3611_149 ),
	.I1(\top/processor/sha_core/n3611_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s128  (
	.I0(\top/processor/sha_core/n3611_153 ),
	.I1(\top/processor/sha_core/n3611_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s129  (
	.I0(\top/processor/sha_core/n3611_157 ),
	.I1(\top/processor/sha_core/n3611_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s130  (
	.I0(\top/processor/sha_core/n3611_161 ),
	.I1(\top/processor/sha_core/n3611_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s131  (
	.I0(\top/processor/sha_core/n3611_133 ),
	.I1(\top/processor/sha_core/n3611_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s132  (
	.I0(\top/processor/sha_core/n3611_137 ),
	.I1(\top/processor/sha_core/n3611_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s133  (
	.I0(\top/processor/sha_core/n3611_141 ),
	.I1(\top/processor/sha_core/n3611_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3709_s134  (
	.I0(\top/processor/sha_core/n3611_145 ),
	.I1(\top/processor/sha_core/n3611_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3709_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s127  (
	.I0(\top/processor/sha_core/n3612_149 ),
	.I1(\top/processor/sha_core/n3612_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s128  (
	.I0(\top/processor/sha_core/n3612_153 ),
	.I1(\top/processor/sha_core/n3612_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s129  (
	.I0(\top/processor/sha_core/n3612_157 ),
	.I1(\top/processor/sha_core/n3612_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s130  (
	.I0(\top/processor/sha_core/n3612_161 ),
	.I1(\top/processor/sha_core/n3612_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s131  (
	.I0(\top/processor/sha_core/n3612_133 ),
	.I1(\top/processor/sha_core/n3612_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s132  (
	.I0(\top/processor/sha_core/n3612_137 ),
	.I1(\top/processor/sha_core/n3612_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s133  (
	.I0(\top/processor/sha_core/n3612_141 ),
	.I1(\top/processor/sha_core/n3612_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3710_s134  (
	.I0(\top/processor/sha_core/n3612_145 ),
	.I1(\top/processor/sha_core/n3612_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3710_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s127  (
	.I0(\top/processor/sha_core/n3613_149 ),
	.I1(\top/processor/sha_core/n3613_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s128  (
	.I0(\top/processor/sha_core/n3613_153 ),
	.I1(\top/processor/sha_core/n3613_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s129  (
	.I0(\top/processor/sha_core/n3613_157 ),
	.I1(\top/processor/sha_core/n3613_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s130  (
	.I0(\top/processor/sha_core/n3613_161 ),
	.I1(\top/processor/sha_core/n3613_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s131  (
	.I0(\top/processor/sha_core/n3613_133 ),
	.I1(\top/processor/sha_core/n3613_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s132  (
	.I0(\top/processor/sha_core/n3613_137 ),
	.I1(\top/processor/sha_core/n3613_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s133  (
	.I0(\top/processor/sha_core/n3613_141 ),
	.I1(\top/processor/sha_core/n3613_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3711_s134  (
	.I0(\top/processor/sha_core/n3613_145 ),
	.I1(\top/processor/sha_core/n3613_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3711_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s127  (
	.I0(\top/processor/sha_core/n3614_149 ),
	.I1(\top/processor/sha_core/n3614_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s128  (
	.I0(\top/processor/sha_core/n3614_153 ),
	.I1(\top/processor/sha_core/n3614_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s129  (
	.I0(\top/processor/sha_core/n3614_157 ),
	.I1(\top/processor/sha_core/n3614_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s130  (
	.I0(\top/processor/sha_core/n3614_161 ),
	.I1(\top/processor/sha_core/n3614_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s131  (
	.I0(\top/processor/sha_core/n3614_133 ),
	.I1(\top/processor/sha_core/n3614_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s132  (
	.I0(\top/processor/sha_core/n3614_137 ),
	.I1(\top/processor/sha_core/n3614_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s133  (
	.I0(\top/processor/sha_core/n3614_141 ),
	.I1(\top/processor/sha_core/n3614_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3712_s134  (
	.I0(\top/processor/sha_core/n3614_145 ),
	.I1(\top/processor/sha_core/n3614_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3712_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s127  (
	.I0(\top/processor/sha_core/n3615_149 ),
	.I1(\top/processor/sha_core/n3615_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s128  (
	.I0(\top/processor/sha_core/n3615_153 ),
	.I1(\top/processor/sha_core/n3615_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s129  (
	.I0(\top/processor/sha_core/n3615_157 ),
	.I1(\top/processor/sha_core/n3615_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s130  (
	.I0(\top/processor/sha_core/n3615_161 ),
	.I1(\top/processor/sha_core/n3615_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s131  (
	.I0(\top/processor/sha_core/n3615_133 ),
	.I1(\top/processor/sha_core/n3615_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s132  (
	.I0(\top/processor/sha_core/n3615_137 ),
	.I1(\top/processor/sha_core/n3615_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s133  (
	.I0(\top/processor/sha_core/n3615_141 ),
	.I1(\top/processor/sha_core/n3615_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3713_s134  (
	.I0(\top/processor/sha_core/n3615_145 ),
	.I1(\top/processor/sha_core/n3615_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3713_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s127  (
	.I0(\top/processor/sha_core/n3616_149 ),
	.I1(\top/processor/sha_core/n3616_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s128  (
	.I0(\top/processor/sha_core/n3616_153 ),
	.I1(\top/processor/sha_core/n3616_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s129  (
	.I0(\top/processor/sha_core/n3616_157 ),
	.I1(\top/processor/sha_core/n3616_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s130  (
	.I0(\top/processor/sha_core/n3616_161 ),
	.I1(\top/processor/sha_core/n3616_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s131  (
	.I0(\top/processor/sha_core/n3616_133 ),
	.I1(\top/processor/sha_core/n3616_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s132  (
	.I0(\top/processor/sha_core/n3616_137 ),
	.I1(\top/processor/sha_core/n3616_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s133  (
	.I0(\top/processor/sha_core/n3616_141 ),
	.I1(\top/processor/sha_core/n3616_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3714_s134  (
	.I0(\top/processor/sha_core/n3616_145 ),
	.I1(\top/processor/sha_core/n3616_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3714_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s127  (
	.I0(\top/processor/sha_core/n3617_149 ),
	.I1(\top/processor/sha_core/n3617_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s128  (
	.I0(\top/processor/sha_core/n3617_153 ),
	.I1(\top/processor/sha_core/n3617_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s129  (
	.I0(\top/processor/sha_core/n3617_157 ),
	.I1(\top/processor/sha_core/n3617_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s130  (
	.I0(\top/processor/sha_core/n3617_161 ),
	.I1(\top/processor/sha_core/n3617_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s131  (
	.I0(\top/processor/sha_core/n3617_133 ),
	.I1(\top/processor/sha_core/n3617_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s132  (
	.I0(\top/processor/sha_core/n3617_137 ),
	.I1(\top/processor/sha_core/n3617_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s133  (
	.I0(\top/processor/sha_core/n3617_141 ),
	.I1(\top/processor/sha_core/n3617_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3715_s134  (
	.I0(\top/processor/sha_core/n3617_145 ),
	.I1(\top/processor/sha_core/n3617_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3715_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s127  (
	.I0(\top/processor/sha_core/n3618_149 ),
	.I1(\top/processor/sha_core/n3618_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s128  (
	.I0(\top/processor/sha_core/n3618_153 ),
	.I1(\top/processor/sha_core/n3618_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s129  (
	.I0(\top/processor/sha_core/n3618_157 ),
	.I1(\top/processor/sha_core/n3618_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s130  (
	.I0(\top/processor/sha_core/n3618_161 ),
	.I1(\top/processor/sha_core/n3618_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s131  (
	.I0(\top/processor/sha_core/n3618_133 ),
	.I1(\top/processor/sha_core/n3618_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s132  (
	.I0(\top/processor/sha_core/n3618_137 ),
	.I1(\top/processor/sha_core/n3618_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s133  (
	.I0(\top/processor/sha_core/n3618_141 ),
	.I1(\top/processor/sha_core/n3618_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3716_s134  (
	.I0(\top/processor/sha_core/n3618_145 ),
	.I1(\top/processor/sha_core/n3618_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3716_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s127  (
	.I0(\top/processor/sha_core/n3619_149 ),
	.I1(\top/processor/sha_core/n3619_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s128  (
	.I0(\top/processor/sha_core/n3619_153 ),
	.I1(\top/processor/sha_core/n3619_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s129  (
	.I0(\top/processor/sha_core/n3619_157 ),
	.I1(\top/processor/sha_core/n3619_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s130  (
	.I0(\top/processor/sha_core/n3619_161 ),
	.I1(\top/processor/sha_core/n3619_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s131  (
	.I0(\top/processor/sha_core/n3619_133 ),
	.I1(\top/processor/sha_core/n3619_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s132  (
	.I0(\top/processor/sha_core/n3619_137 ),
	.I1(\top/processor/sha_core/n3619_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s133  (
	.I0(\top/processor/sha_core/n3619_141 ),
	.I1(\top/processor/sha_core/n3619_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3717_s134  (
	.I0(\top/processor/sha_core/n3619_145 ),
	.I1(\top/processor/sha_core/n3619_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3717_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s127  (
	.I0(\top/processor/sha_core/n3620_149 ),
	.I1(\top/processor/sha_core/n3620_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s128  (
	.I0(\top/processor/sha_core/n3620_153 ),
	.I1(\top/processor/sha_core/n3620_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s129  (
	.I0(\top/processor/sha_core/n3620_157 ),
	.I1(\top/processor/sha_core/n3620_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s130  (
	.I0(\top/processor/sha_core/n3620_161 ),
	.I1(\top/processor/sha_core/n3620_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s131  (
	.I0(\top/processor/sha_core/n3620_133 ),
	.I1(\top/processor/sha_core/n3620_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s132  (
	.I0(\top/processor/sha_core/n3620_137 ),
	.I1(\top/processor/sha_core/n3620_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s133  (
	.I0(\top/processor/sha_core/n3620_141 ),
	.I1(\top/processor/sha_core/n3620_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3718_s134  (
	.I0(\top/processor/sha_core/n3620_145 ),
	.I1(\top/processor/sha_core/n3620_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3718_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s127  (
	.I0(\top/processor/sha_core/n3621_149 ),
	.I1(\top/processor/sha_core/n3621_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s128  (
	.I0(\top/processor/sha_core/n3621_153 ),
	.I1(\top/processor/sha_core/n3621_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s129  (
	.I0(\top/processor/sha_core/n3621_157 ),
	.I1(\top/processor/sha_core/n3621_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s130  (
	.I0(\top/processor/sha_core/n3621_161 ),
	.I1(\top/processor/sha_core/n3621_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s131  (
	.I0(\top/processor/sha_core/n3621_133 ),
	.I1(\top/processor/sha_core/n3621_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s132  (
	.I0(\top/processor/sha_core/n3621_137 ),
	.I1(\top/processor/sha_core/n3621_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s133  (
	.I0(\top/processor/sha_core/n3621_141 ),
	.I1(\top/processor/sha_core/n3621_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3719_s134  (
	.I0(\top/processor/sha_core/n3621_145 ),
	.I1(\top/processor/sha_core/n3621_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3719_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s127  (
	.I0(\top/processor/sha_core/n3622_149 ),
	.I1(\top/processor/sha_core/n3622_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s128  (
	.I0(\top/processor/sha_core/n3622_153 ),
	.I1(\top/processor/sha_core/n3622_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s129  (
	.I0(\top/processor/sha_core/n3622_157 ),
	.I1(\top/processor/sha_core/n3622_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s130  (
	.I0(\top/processor/sha_core/n3622_161 ),
	.I1(\top/processor/sha_core/n3622_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s131  (
	.I0(\top/processor/sha_core/n3622_133 ),
	.I1(\top/processor/sha_core/n3622_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s132  (
	.I0(\top/processor/sha_core/n3622_137 ),
	.I1(\top/processor/sha_core/n3622_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s133  (
	.I0(\top/processor/sha_core/n3622_141 ),
	.I1(\top/processor/sha_core/n3622_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3720_s134  (
	.I0(\top/processor/sha_core/n3622_145 ),
	.I1(\top/processor/sha_core/n3622_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3720_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s127  (
	.I0(\top/processor/sha_core/n3623_149 ),
	.I1(\top/processor/sha_core/n3623_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s128  (
	.I0(\top/processor/sha_core/n3623_153 ),
	.I1(\top/processor/sha_core/n3623_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s129  (
	.I0(\top/processor/sha_core/n3623_157 ),
	.I1(\top/processor/sha_core/n3623_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s130  (
	.I0(\top/processor/sha_core/n3623_161 ),
	.I1(\top/processor/sha_core/n3623_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s131  (
	.I0(\top/processor/sha_core/n3623_133 ),
	.I1(\top/processor/sha_core/n3623_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s132  (
	.I0(\top/processor/sha_core/n3623_137 ),
	.I1(\top/processor/sha_core/n3623_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s133  (
	.I0(\top/processor/sha_core/n3623_141 ),
	.I1(\top/processor/sha_core/n3623_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3721_s134  (
	.I0(\top/processor/sha_core/n3623_145 ),
	.I1(\top/processor/sha_core/n3623_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3721_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s127  (
	.I0(\top/processor/sha_core/n3624_149 ),
	.I1(\top/processor/sha_core/n3624_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s128  (
	.I0(\top/processor/sha_core/n3624_153 ),
	.I1(\top/processor/sha_core/n3624_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s129  (
	.I0(\top/processor/sha_core/n3624_157 ),
	.I1(\top/processor/sha_core/n3624_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s130  (
	.I0(\top/processor/sha_core/n3624_161 ),
	.I1(\top/processor/sha_core/n3624_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s131  (
	.I0(\top/processor/sha_core/n3624_133 ),
	.I1(\top/processor/sha_core/n3624_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s132  (
	.I0(\top/processor/sha_core/n3624_137 ),
	.I1(\top/processor/sha_core/n3624_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s133  (
	.I0(\top/processor/sha_core/n3624_141 ),
	.I1(\top/processor/sha_core/n3624_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3722_s134  (
	.I0(\top/processor/sha_core/n3624_145 ),
	.I1(\top/processor/sha_core/n3624_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3722_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s127  (
	.I0(\top/processor/sha_core/n3625_149 ),
	.I1(\top/processor/sha_core/n3625_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s128  (
	.I0(\top/processor/sha_core/n3625_153 ),
	.I1(\top/processor/sha_core/n3625_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s129  (
	.I0(\top/processor/sha_core/n3625_157 ),
	.I1(\top/processor/sha_core/n3625_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s130  (
	.I0(\top/processor/sha_core/n3625_161 ),
	.I1(\top/processor/sha_core/n3625_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s131  (
	.I0(\top/processor/sha_core/n3625_133 ),
	.I1(\top/processor/sha_core/n3625_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s132  (
	.I0(\top/processor/sha_core/n3625_137 ),
	.I1(\top/processor/sha_core/n3625_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s133  (
	.I0(\top/processor/sha_core/n3625_141 ),
	.I1(\top/processor/sha_core/n3625_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3723_s134  (
	.I0(\top/processor/sha_core/n3625_145 ),
	.I1(\top/processor/sha_core/n3625_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3723_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s127  (
	.I0(\top/processor/sha_core/n3626_149 ),
	.I1(\top/processor/sha_core/n3626_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s128  (
	.I0(\top/processor/sha_core/n3626_153 ),
	.I1(\top/processor/sha_core/n3626_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s129  (
	.I0(\top/processor/sha_core/n3626_157 ),
	.I1(\top/processor/sha_core/n3626_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s130  (
	.I0(\top/processor/sha_core/n3626_161 ),
	.I1(\top/processor/sha_core/n3626_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s131  (
	.I0(\top/processor/sha_core/n3626_133 ),
	.I1(\top/processor/sha_core/n3626_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s132  (
	.I0(\top/processor/sha_core/n3626_137 ),
	.I1(\top/processor/sha_core/n3626_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s133  (
	.I0(\top/processor/sha_core/n3626_141 ),
	.I1(\top/processor/sha_core/n3626_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3724_s134  (
	.I0(\top/processor/sha_core/n3626_145 ),
	.I1(\top/processor/sha_core/n3626_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3724_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s127  (
	.I0(\top/processor/sha_core/n3627_149 ),
	.I1(\top/processor/sha_core/n3627_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s128  (
	.I0(\top/processor/sha_core/n3627_153 ),
	.I1(\top/processor/sha_core/n3627_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s129  (
	.I0(\top/processor/sha_core/n3627_157 ),
	.I1(\top/processor/sha_core/n3627_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s130  (
	.I0(\top/processor/sha_core/n3627_161 ),
	.I1(\top/processor/sha_core/n3627_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s131  (
	.I0(\top/processor/sha_core/n3627_133 ),
	.I1(\top/processor/sha_core/n3627_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s132  (
	.I0(\top/processor/sha_core/n3627_137 ),
	.I1(\top/processor/sha_core/n3627_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s133  (
	.I0(\top/processor/sha_core/n3627_141 ),
	.I1(\top/processor/sha_core/n3627_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3725_s134  (
	.I0(\top/processor/sha_core/n3627_145 ),
	.I1(\top/processor/sha_core/n3627_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3725_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s127  (
	.I0(\top/processor/sha_core/n3628_149 ),
	.I1(\top/processor/sha_core/n3628_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s128  (
	.I0(\top/processor/sha_core/n3628_153 ),
	.I1(\top/processor/sha_core/n3628_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s129  (
	.I0(\top/processor/sha_core/n3628_157 ),
	.I1(\top/processor/sha_core/n3628_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s130  (
	.I0(\top/processor/sha_core/n3628_161 ),
	.I1(\top/processor/sha_core/n3628_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s131  (
	.I0(\top/processor/sha_core/n3628_133 ),
	.I1(\top/processor/sha_core/n3628_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s132  (
	.I0(\top/processor/sha_core/n3628_137 ),
	.I1(\top/processor/sha_core/n3628_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s133  (
	.I0(\top/processor/sha_core/n3628_141 ),
	.I1(\top/processor/sha_core/n3628_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3726_s134  (
	.I0(\top/processor/sha_core/n3628_145 ),
	.I1(\top/processor/sha_core/n3628_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3726_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s127  (
	.I0(\top/processor/sha_core/n3629_149 ),
	.I1(\top/processor/sha_core/n3629_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s128  (
	.I0(\top/processor/sha_core/n3629_153 ),
	.I1(\top/processor/sha_core/n3629_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s129  (
	.I0(\top/processor/sha_core/n3629_157 ),
	.I1(\top/processor/sha_core/n3629_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s130  (
	.I0(\top/processor/sha_core/n3629_161 ),
	.I1(\top/processor/sha_core/n3629_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s131  (
	.I0(\top/processor/sha_core/n3629_133 ),
	.I1(\top/processor/sha_core/n3629_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s132  (
	.I0(\top/processor/sha_core/n3629_137 ),
	.I1(\top/processor/sha_core/n3629_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s133  (
	.I0(\top/processor/sha_core/n3629_141 ),
	.I1(\top/processor/sha_core/n3629_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3727_s134  (
	.I0(\top/processor/sha_core/n3629_145 ),
	.I1(\top/processor/sha_core/n3629_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3727_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s127  (
	.I0(\top/processor/sha_core/n3630_149 ),
	.I1(\top/processor/sha_core/n3630_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s128  (
	.I0(\top/processor/sha_core/n3630_153 ),
	.I1(\top/processor/sha_core/n3630_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s129  (
	.I0(\top/processor/sha_core/n3630_157 ),
	.I1(\top/processor/sha_core/n3630_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s130  (
	.I0(\top/processor/sha_core/n3630_161 ),
	.I1(\top/processor/sha_core/n3630_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s131  (
	.I0(\top/processor/sha_core/n3630_133 ),
	.I1(\top/processor/sha_core/n3630_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s132  (
	.I0(\top/processor/sha_core/n3630_137 ),
	.I1(\top/processor/sha_core/n3630_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s133  (
	.I0(\top/processor/sha_core/n3630_141 ),
	.I1(\top/processor/sha_core/n3630_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3728_s134  (
	.I0(\top/processor/sha_core/n3630_145 ),
	.I1(\top/processor/sha_core/n3630_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3728_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s127  (
	.I0(\top/processor/sha_core/n3631_149 ),
	.I1(\top/processor/sha_core/n3631_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s128  (
	.I0(\top/processor/sha_core/n3631_153 ),
	.I1(\top/processor/sha_core/n3631_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s129  (
	.I0(\top/processor/sha_core/n3631_157 ),
	.I1(\top/processor/sha_core/n3631_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s130  (
	.I0(\top/processor/sha_core/n3631_161 ),
	.I1(\top/processor/sha_core/n3631_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s131  (
	.I0(\top/processor/sha_core/n3631_133 ),
	.I1(\top/processor/sha_core/n3631_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s132  (
	.I0(\top/processor/sha_core/n3631_137 ),
	.I1(\top/processor/sha_core/n3631_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s133  (
	.I0(\top/processor/sha_core/n3631_141 ),
	.I1(\top/processor/sha_core/n3631_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3729_s134  (
	.I0(\top/processor/sha_core/n3631_145 ),
	.I1(\top/processor/sha_core/n3631_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3729_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s127  (
	.I0(\top/processor/sha_core/n3632_149 ),
	.I1(\top/processor/sha_core/n3632_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s128  (
	.I0(\top/processor/sha_core/n3632_153 ),
	.I1(\top/processor/sha_core/n3632_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s129  (
	.I0(\top/processor/sha_core/n3632_157 ),
	.I1(\top/processor/sha_core/n3632_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s130  (
	.I0(\top/processor/sha_core/n3632_161 ),
	.I1(\top/processor/sha_core/n3632_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s131  (
	.I0(\top/processor/sha_core/n3632_133 ),
	.I1(\top/processor/sha_core/n3632_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s132  (
	.I0(\top/processor/sha_core/n3632_137 ),
	.I1(\top/processor/sha_core/n3632_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s133  (
	.I0(\top/processor/sha_core/n3632_141 ),
	.I1(\top/processor/sha_core/n3632_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3730_s134  (
	.I0(\top/processor/sha_core/n3632_145 ),
	.I1(\top/processor/sha_core/n3632_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3730_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s127  (
	.I0(\top/processor/sha_core/n3633_149 ),
	.I1(\top/processor/sha_core/n3633_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s128  (
	.I0(\top/processor/sha_core/n3633_153 ),
	.I1(\top/processor/sha_core/n3633_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s129  (
	.I0(\top/processor/sha_core/n3633_157 ),
	.I1(\top/processor/sha_core/n3633_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s130  (
	.I0(\top/processor/sha_core/n3633_161 ),
	.I1(\top/processor/sha_core/n3633_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s131  (
	.I0(\top/processor/sha_core/n3633_133 ),
	.I1(\top/processor/sha_core/n3633_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s132  (
	.I0(\top/processor/sha_core/n3633_137 ),
	.I1(\top/processor/sha_core/n3633_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s133  (
	.I0(\top/processor/sha_core/n3633_141 ),
	.I1(\top/processor/sha_core/n3633_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3731_s134  (
	.I0(\top/processor/sha_core/n3633_145 ),
	.I1(\top/processor/sha_core/n3633_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3731_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s127  (
	.I0(\top/processor/sha_core/n3634_149 ),
	.I1(\top/processor/sha_core/n3634_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s128  (
	.I0(\top/processor/sha_core/n3634_153 ),
	.I1(\top/processor/sha_core/n3634_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s129  (
	.I0(\top/processor/sha_core/n3634_157 ),
	.I1(\top/processor/sha_core/n3634_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s130  (
	.I0(\top/processor/sha_core/n3634_161 ),
	.I1(\top/processor/sha_core/n3634_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s131  (
	.I0(\top/processor/sha_core/n3634_133 ),
	.I1(\top/processor/sha_core/n3634_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s132  (
	.I0(\top/processor/sha_core/n3634_137 ),
	.I1(\top/processor/sha_core/n3634_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s133  (
	.I0(\top/processor/sha_core/n3634_141 ),
	.I1(\top/processor/sha_core/n3634_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3732_s134  (
	.I0(\top/processor/sha_core/n3634_145 ),
	.I1(\top/processor/sha_core/n3634_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3732_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s127  (
	.I0(\top/processor/sha_core/n3635_149 ),
	.I1(\top/processor/sha_core/n3635_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s128  (
	.I0(\top/processor/sha_core/n3635_153 ),
	.I1(\top/processor/sha_core/n3635_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s129  (
	.I0(\top/processor/sha_core/n3635_157 ),
	.I1(\top/processor/sha_core/n3635_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s130  (
	.I0(\top/processor/sha_core/n3635_161 ),
	.I1(\top/processor/sha_core/n3635_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s131  (
	.I0(\top/processor/sha_core/n3635_133 ),
	.I1(\top/processor/sha_core/n3635_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s132  (
	.I0(\top/processor/sha_core/n3635_137 ),
	.I1(\top/processor/sha_core/n3635_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s133  (
	.I0(\top/processor/sha_core/n3635_141 ),
	.I1(\top/processor/sha_core/n3635_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3733_s134  (
	.I0(\top/processor/sha_core/n3635_145 ),
	.I1(\top/processor/sha_core/n3635_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3733_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s127  (
	.I0(\top/processor/sha_core/n3636_149 ),
	.I1(\top/processor/sha_core/n3636_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s128  (
	.I0(\top/processor/sha_core/n3636_153 ),
	.I1(\top/processor/sha_core/n3636_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s129  (
	.I0(\top/processor/sha_core/n3636_157 ),
	.I1(\top/processor/sha_core/n3636_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s130  (
	.I0(\top/processor/sha_core/n3636_161 ),
	.I1(\top/processor/sha_core/n3636_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s131  (
	.I0(\top/processor/sha_core/n3636_133 ),
	.I1(\top/processor/sha_core/n3636_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s132  (
	.I0(\top/processor/sha_core/n3636_137 ),
	.I1(\top/processor/sha_core/n3636_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s133  (
	.I0(\top/processor/sha_core/n3636_141 ),
	.I1(\top/processor/sha_core/n3636_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3734_s134  (
	.I0(\top/processor/sha_core/n3636_145 ),
	.I1(\top/processor/sha_core/n3636_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3734_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s127  (
	.I0(\top/processor/sha_core/n3637_149 ),
	.I1(\top/processor/sha_core/n3637_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s128  (
	.I0(\top/processor/sha_core/n3637_153 ),
	.I1(\top/processor/sha_core/n3637_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s129  (
	.I0(\top/processor/sha_core/n3637_157 ),
	.I1(\top/processor/sha_core/n3637_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s130  (
	.I0(\top/processor/sha_core/n3637_161 ),
	.I1(\top/processor/sha_core/n3637_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s131  (
	.I0(\top/processor/sha_core/n3637_133 ),
	.I1(\top/processor/sha_core/n3637_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s132  (
	.I0(\top/processor/sha_core/n3637_137 ),
	.I1(\top/processor/sha_core/n3637_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s133  (
	.I0(\top/processor/sha_core/n3637_141 ),
	.I1(\top/processor/sha_core/n3637_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3735_s134  (
	.I0(\top/processor/sha_core/n3637_145 ),
	.I1(\top/processor/sha_core/n3637_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3735_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s127  (
	.I0(\top/processor/sha_core/n3638_149 ),
	.I1(\top/processor/sha_core/n3638_151 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s128  (
	.I0(\top/processor/sha_core/n3638_153 ),
	.I1(\top/processor/sha_core/n3638_155 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s129  (
	.I0(\top/processor/sha_core/n3638_157 ),
	.I1(\top/processor/sha_core/n3638_159 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s130  (
	.I0(\top/processor/sha_core/n3638_161 ),
	.I1(\top/processor/sha_core/n3638_163 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s131  (
	.I0(\top/processor/sha_core/n3638_133 ),
	.I1(\top/processor/sha_core/n3638_135 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_141 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s132  (
	.I0(\top/processor/sha_core/n3638_137 ),
	.I1(\top/processor/sha_core/n3638_139 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_143 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s133  (
	.I0(\top/processor/sha_core/n3638_141 ),
	.I1(\top/processor/sha_core/n3638_143 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_145 )
);
MUX2_LUT5 \top/processor/sha_core/n3736_s134  (
	.I0(\top/processor/sha_core/n3638_145 ),
	.I1(\top/processor/sha_core/n3638_147 ),
	.S0(\top/processor/sha_core/n3452_7 ),
	.O(\top/processor/sha_core/n3736_147 )
);
MUX2_LUT5 \top/processor/sha_core/n3860_s129  (
	.I0(\top/processor/sha_core/n3860_107 ),
	.I1(\top/processor/sha_core/n3860_109 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3860_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3860_s128  (
	.I0(\top/processor/sha_core/n3860_111 ),
	.I1(\top/processor/sha_core/n3860_113 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3860_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3860_s131  (
	.I0(\top/processor/sha_core/n3860_115 ),
	.I1(\top/processor/sha_core/n3860_101 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3860_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3860_s130  (
	.I0(\top/processor/sha_core/n3860_103 ),
	.I1(\top/processor/sha_core/n3860_105 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3860_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3861_s129  (
	.I0(\top/processor/sha_core/n3861_101 ),
	.I1(\top/processor/sha_core/n3861_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3861_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3861_s128  (
	.I0(\top/processor/sha_core/n3861_105 ),
	.I1(\top/processor/sha_core/n3861_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3861_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3861_s131  (
	.I0(\top/processor/sha_core/n3861_109 ),
	.I1(\top/processor/sha_core/n3861_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3861_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3861_s130  (
	.I0(\top/processor/sha_core/n3861_113 ),
	.I1(\top/processor/sha_core/n3861_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3861_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3862_s129  (
	.I0(\top/processor/sha_core/n3862_101 ),
	.I1(\top/processor/sha_core/n3862_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3862_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3862_s128  (
	.I0(\top/processor/sha_core/n3862_105 ),
	.I1(\top/processor/sha_core/n3862_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3862_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3862_s131  (
	.I0(\top/processor/sha_core/n3862_109 ),
	.I1(\top/processor/sha_core/n3862_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3862_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3862_s130  (
	.I0(\top/processor/sha_core/n3862_113 ),
	.I1(\top/processor/sha_core/n3862_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3862_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3863_s129  (
	.I0(\top/processor/sha_core/n3863_101 ),
	.I1(\top/processor/sha_core/n3863_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3863_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3863_s128  (
	.I0(\top/processor/sha_core/n3863_105 ),
	.I1(\top/processor/sha_core/n3863_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3863_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3863_s131  (
	.I0(\top/processor/sha_core/n3863_109 ),
	.I1(\top/processor/sha_core/n3863_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3863_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3863_s130  (
	.I0(\top/processor/sha_core/n3863_113 ),
	.I1(\top/processor/sha_core/n3863_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3863_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3864_s129  (
	.I0(\top/processor/sha_core/n3864_101 ),
	.I1(\top/processor/sha_core/n3864_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3864_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3864_s128  (
	.I0(\top/processor/sha_core/n3864_105 ),
	.I1(\top/processor/sha_core/n3864_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3864_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3864_s131  (
	.I0(\top/processor/sha_core/n3864_109 ),
	.I1(\top/processor/sha_core/n3864_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3864_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3864_s130  (
	.I0(\top/processor/sha_core/n3864_113 ),
	.I1(\top/processor/sha_core/n3864_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3864_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3865_s129  (
	.I0(\top/processor/sha_core/n3865_101 ),
	.I1(\top/processor/sha_core/n3865_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3865_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3865_s128  (
	.I0(\top/processor/sha_core/n3865_105 ),
	.I1(\top/processor/sha_core/n3865_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3865_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3865_s131  (
	.I0(\top/processor/sha_core/n3865_109 ),
	.I1(\top/processor/sha_core/n3865_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3865_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3865_s130  (
	.I0(\top/processor/sha_core/n3865_113 ),
	.I1(\top/processor/sha_core/n3865_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3865_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3866_s129  (
	.I0(\top/processor/sha_core/n3866_113 ),
	.I1(\top/processor/sha_core/n3866_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3866_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3866_s128  (
	.I0(\top/processor/sha_core/n3866_101 ),
	.I1(\top/processor/sha_core/n3866_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3866_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3866_s131  (
	.I0(\top/processor/sha_core/n3866_105 ),
	.I1(\top/processor/sha_core/n3866_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3866_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3866_s130  (
	.I0(\top/processor/sha_core/n3866_109 ),
	.I1(\top/processor/sha_core/n3866_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3866_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3867_s129  (
	.I0(\top/processor/sha_core/n3867_101 ),
	.I1(\top/processor/sha_core/n3867_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3867_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3867_s128  (
	.I0(\top/processor/sha_core/n3867_105 ),
	.I1(\top/processor/sha_core/n3867_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3867_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3867_s131  (
	.I0(\top/processor/sha_core/n3867_109 ),
	.I1(\top/processor/sha_core/n3867_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3867_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3867_s130  (
	.I0(\top/processor/sha_core/n3867_113 ),
	.I1(\top/processor/sha_core/n3867_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3867_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3868_s129  (
	.I0(\top/processor/sha_core/n3868_101 ),
	.I1(\top/processor/sha_core/n3868_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3868_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3868_s128  (
	.I0(\top/processor/sha_core/n3868_105 ),
	.I1(\top/processor/sha_core/n3868_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3868_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3868_s131  (
	.I0(\top/processor/sha_core/n3868_109 ),
	.I1(\top/processor/sha_core/n3868_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3868_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3868_s130  (
	.I0(\top/processor/sha_core/n3868_113 ),
	.I1(\top/processor/sha_core/n3868_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3868_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3869_s129  (
	.I0(\top/processor/sha_core/n3869_101 ),
	.I1(\top/processor/sha_core/n3869_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3869_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3869_s128  (
	.I0(\top/processor/sha_core/n3869_105 ),
	.I1(\top/processor/sha_core/n3869_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3869_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3869_s131  (
	.I0(\top/processor/sha_core/n3869_109 ),
	.I1(\top/processor/sha_core/n3869_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3869_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3869_s130  (
	.I0(\top/processor/sha_core/n3869_113 ),
	.I1(\top/processor/sha_core/n3869_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3869_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3870_s129  (
	.I0(\top/processor/sha_core/n3870_101 ),
	.I1(\top/processor/sha_core/n3870_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3870_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3870_s128  (
	.I0(\top/processor/sha_core/n3870_105 ),
	.I1(\top/processor/sha_core/n3870_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3870_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3870_s131  (
	.I0(\top/processor/sha_core/n3870_109 ),
	.I1(\top/processor/sha_core/n3870_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3870_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3870_s130  (
	.I0(\top/processor/sha_core/n3870_113 ),
	.I1(\top/processor/sha_core/n3870_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3870_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3871_s129  (
	.I0(\top/processor/sha_core/n3871_101 ),
	.I1(\top/processor/sha_core/n3871_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3871_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3871_s128  (
	.I0(\top/processor/sha_core/n3871_105 ),
	.I1(\top/processor/sha_core/n3871_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3871_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3871_s131  (
	.I0(\top/processor/sha_core/n3871_109 ),
	.I1(\top/processor/sha_core/n3871_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3871_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3871_s130  (
	.I0(\top/processor/sha_core/n3871_113 ),
	.I1(\top/processor/sha_core/n3871_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3871_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3872_s129  (
	.I0(\top/processor/sha_core/n3872_101 ),
	.I1(\top/processor/sha_core/n3872_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3872_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3872_s128  (
	.I0(\top/processor/sha_core/n3872_105 ),
	.I1(\top/processor/sha_core/n3872_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3872_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3872_s131  (
	.I0(\top/processor/sha_core/n3872_109 ),
	.I1(\top/processor/sha_core/n3872_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3872_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3872_s130  (
	.I0(\top/processor/sha_core/n3872_113 ),
	.I1(\top/processor/sha_core/n3872_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3872_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3873_s129  (
	.I0(\top/processor/sha_core/n3873_101 ),
	.I1(\top/processor/sha_core/n3873_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3873_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3873_s128  (
	.I0(\top/processor/sha_core/n3873_105 ),
	.I1(\top/processor/sha_core/n3873_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3873_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3873_s131  (
	.I0(\top/processor/sha_core/n3873_109 ),
	.I1(\top/processor/sha_core/n3873_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3873_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3873_s130  (
	.I0(\top/processor/sha_core/n3873_113 ),
	.I1(\top/processor/sha_core/n3873_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3873_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3874_s129  (
	.I0(\top/processor/sha_core/n3874_101 ),
	.I1(\top/processor/sha_core/n3874_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3874_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3874_s128  (
	.I0(\top/processor/sha_core/n3874_105 ),
	.I1(\top/processor/sha_core/n3874_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3874_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3874_s131  (
	.I0(\top/processor/sha_core/n3874_109 ),
	.I1(\top/processor/sha_core/n3874_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3874_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3874_s130  (
	.I0(\top/processor/sha_core/n3874_113 ),
	.I1(\top/processor/sha_core/n3874_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3874_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3875_s129  (
	.I0(\top/processor/sha_core/n3875_101 ),
	.I1(\top/processor/sha_core/n3875_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3875_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3875_s128  (
	.I0(\top/processor/sha_core/n3875_105 ),
	.I1(\top/processor/sha_core/n3875_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3875_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3875_s131  (
	.I0(\top/processor/sha_core/n3875_109 ),
	.I1(\top/processor/sha_core/n3875_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3875_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3875_s130  (
	.I0(\top/processor/sha_core/n3875_113 ),
	.I1(\top/processor/sha_core/n3875_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3875_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3876_s129  (
	.I0(\top/processor/sha_core/n3876_101 ),
	.I1(\top/processor/sha_core/n3876_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3876_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3876_s128  (
	.I0(\top/processor/sha_core/n3876_105 ),
	.I1(\top/processor/sha_core/n3876_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3876_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3876_s131  (
	.I0(\top/processor/sha_core/n3876_109 ),
	.I1(\top/processor/sha_core/n3876_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3876_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3876_s130  (
	.I0(\top/processor/sha_core/n3876_113 ),
	.I1(\top/processor/sha_core/n3876_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3876_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3877_s129  (
	.I0(\top/processor/sha_core/n3877_101 ),
	.I1(\top/processor/sha_core/n3877_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3877_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3877_s128  (
	.I0(\top/processor/sha_core/n3877_105 ),
	.I1(\top/processor/sha_core/n3877_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3877_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3877_s131  (
	.I0(\top/processor/sha_core/n3877_109 ),
	.I1(\top/processor/sha_core/n3877_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3877_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3877_s130  (
	.I0(\top/processor/sha_core/n3877_113 ),
	.I1(\top/processor/sha_core/n3877_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3877_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3878_s129  (
	.I0(\top/processor/sha_core/n3878_101 ),
	.I1(\top/processor/sha_core/n3878_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3878_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3878_s128  (
	.I0(\top/processor/sha_core/n3878_105 ),
	.I1(\top/processor/sha_core/n3878_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3878_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3878_s131  (
	.I0(\top/processor/sha_core/n3878_109 ),
	.I1(\top/processor/sha_core/n3878_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3878_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3878_s130  (
	.I0(\top/processor/sha_core/n3878_113 ),
	.I1(\top/processor/sha_core/n3878_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3878_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3879_s129  (
	.I0(\top/processor/sha_core/n3879_101 ),
	.I1(\top/processor/sha_core/n3879_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3879_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3879_s128  (
	.I0(\top/processor/sha_core/n3879_105 ),
	.I1(\top/processor/sha_core/n3879_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3879_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3879_s131  (
	.I0(\top/processor/sha_core/n3879_109 ),
	.I1(\top/processor/sha_core/n3879_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3879_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3879_s130  (
	.I0(\top/processor/sha_core/n3879_113 ),
	.I1(\top/processor/sha_core/n3879_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3879_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3880_s129  (
	.I0(\top/processor/sha_core/n3880_101 ),
	.I1(\top/processor/sha_core/n3880_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3880_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3880_s128  (
	.I0(\top/processor/sha_core/n3880_105 ),
	.I1(\top/processor/sha_core/n3880_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3880_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3880_s131  (
	.I0(\top/processor/sha_core/n3880_109 ),
	.I1(\top/processor/sha_core/n3880_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3880_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3880_s130  (
	.I0(\top/processor/sha_core/n3880_113 ),
	.I1(\top/processor/sha_core/n3880_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3880_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3881_s129  (
	.I0(\top/processor/sha_core/n3881_101 ),
	.I1(\top/processor/sha_core/n3881_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3881_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3881_s128  (
	.I0(\top/processor/sha_core/n3881_105 ),
	.I1(\top/processor/sha_core/n3881_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3881_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3881_s131  (
	.I0(\top/processor/sha_core/n3881_109 ),
	.I1(\top/processor/sha_core/n3881_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3881_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3881_s130  (
	.I0(\top/processor/sha_core/n3881_113 ),
	.I1(\top/processor/sha_core/n3881_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3881_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3882_s129  (
	.I0(\top/processor/sha_core/n3882_101 ),
	.I1(\top/processor/sha_core/n3882_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3882_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3882_s128  (
	.I0(\top/processor/sha_core/n3882_105 ),
	.I1(\top/processor/sha_core/n3882_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3882_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3882_s131  (
	.I0(\top/processor/sha_core/n3882_109 ),
	.I1(\top/processor/sha_core/n3882_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3882_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3882_s130  (
	.I0(\top/processor/sha_core/n3882_113 ),
	.I1(\top/processor/sha_core/n3882_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3882_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3883_s129  (
	.I0(\top/processor/sha_core/n3883_101 ),
	.I1(\top/processor/sha_core/n3883_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3883_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3883_s128  (
	.I0(\top/processor/sha_core/n3883_105 ),
	.I1(\top/processor/sha_core/n3883_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3883_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3883_s131  (
	.I0(\top/processor/sha_core/n3883_109 ),
	.I1(\top/processor/sha_core/n3883_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3883_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3883_s130  (
	.I0(\top/processor/sha_core/n3883_113 ),
	.I1(\top/processor/sha_core/n3883_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3883_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3884_s129  (
	.I0(\top/processor/sha_core/n3884_101 ),
	.I1(\top/processor/sha_core/n3884_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3884_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3884_s128  (
	.I0(\top/processor/sha_core/n3884_105 ),
	.I1(\top/processor/sha_core/n3884_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3884_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3884_s131  (
	.I0(\top/processor/sha_core/n3884_109 ),
	.I1(\top/processor/sha_core/n3884_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3884_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3884_s130  (
	.I0(\top/processor/sha_core/n3884_113 ),
	.I1(\top/processor/sha_core/n3884_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3884_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3885_s129  (
	.I0(\top/processor/sha_core/n3885_101 ),
	.I1(\top/processor/sha_core/n3885_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3885_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3885_s128  (
	.I0(\top/processor/sha_core/n3885_105 ),
	.I1(\top/processor/sha_core/n3885_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3885_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3885_s131  (
	.I0(\top/processor/sha_core/n3885_109 ),
	.I1(\top/processor/sha_core/n3885_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3885_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3885_s130  (
	.I0(\top/processor/sha_core/n3885_113 ),
	.I1(\top/processor/sha_core/n3885_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3885_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3886_s129  (
	.I0(\top/processor/sha_core/n3886_101 ),
	.I1(\top/processor/sha_core/n3886_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3886_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3886_s128  (
	.I0(\top/processor/sha_core/n3886_105 ),
	.I1(\top/processor/sha_core/n3886_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3886_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3886_s131  (
	.I0(\top/processor/sha_core/n3886_109 ),
	.I1(\top/processor/sha_core/n3886_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3886_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3886_s130  (
	.I0(\top/processor/sha_core/n3886_113 ),
	.I1(\top/processor/sha_core/n3886_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3886_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3887_s129  (
	.I0(\top/processor/sha_core/n3887_101 ),
	.I1(\top/processor/sha_core/n3887_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3887_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3887_s128  (
	.I0(\top/processor/sha_core/n3887_105 ),
	.I1(\top/processor/sha_core/n3887_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3887_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3887_s131  (
	.I0(\top/processor/sha_core/n3887_109 ),
	.I1(\top/processor/sha_core/n3887_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3887_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3887_s130  (
	.I0(\top/processor/sha_core/n3887_113 ),
	.I1(\top/processor/sha_core/n3887_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3887_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3888_s129  (
	.I0(\top/processor/sha_core/n3888_101 ),
	.I1(\top/processor/sha_core/n3888_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3888_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3888_s128  (
	.I0(\top/processor/sha_core/n3888_105 ),
	.I1(\top/processor/sha_core/n3888_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3888_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3888_s131  (
	.I0(\top/processor/sha_core/n3888_109 ),
	.I1(\top/processor/sha_core/n3888_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3888_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3888_s130  (
	.I0(\top/processor/sha_core/n3888_113 ),
	.I1(\top/processor/sha_core/n3888_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3888_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3889_s129  (
	.I0(\top/processor/sha_core/n3889_101 ),
	.I1(\top/processor/sha_core/n3889_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3889_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3889_s128  (
	.I0(\top/processor/sha_core/n3889_105 ),
	.I1(\top/processor/sha_core/n3889_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3889_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3889_s131  (
	.I0(\top/processor/sha_core/n3889_109 ),
	.I1(\top/processor/sha_core/n3889_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3889_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3889_s130  (
	.I0(\top/processor/sha_core/n3889_113 ),
	.I1(\top/processor/sha_core/n3889_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3889_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3890_s129  (
	.I0(\top/processor/sha_core/n3890_101 ),
	.I1(\top/processor/sha_core/n3890_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3890_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3890_s128  (
	.I0(\top/processor/sha_core/n3890_105 ),
	.I1(\top/processor/sha_core/n3890_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3890_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3890_s131  (
	.I0(\top/processor/sha_core/n3890_109 ),
	.I1(\top/processor/sha_core/n3890_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3890_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3890_s130  (
	.I0(\top/processor/sha_core/n3890_113 ),
	.I1(\top/processor/sha_core/n3890_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3890_139 )
);
MUX2_LUT5 \top/processor/sha_core/n3891_s129  (
	.I0(\top/processor/sha_core/n3891_101 ),
	.I1(\top/processor/sha_core/n3891_103 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3891_133 )
);
MUX2_LUT5 \top/processor/sha_core/n3891_s128  (
	.I0(\top/processor/sha_core/n3891_105 ),
	.I1(\top/processor/sha_core/n3891_107 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3891_135 )
);
MUX2_LUT5 \top/processor/sha_core/n3891_s131  (
	.I0(\top/processor/sha_core/n3891_109 ),
	.I1(\top/processor/sha_core/n3891_111 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3891_137 )
);
MUX2_LUT5 \top/processor/sha_core/n3891_s130  (
	.I0(\top/processor/sha_core/n3891_113 ),
	.I1(\top/processor/sha_core/n3891_115 ),
	.S0(\top/processor/sha_core/msg_idx [3]),
	.O(\top/processor/sha_core/n3891_139 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s194  (
	.I0(\top/processor/sha_core/n327_165 ),
	.I1(\top/processor/sha_core/n327_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_197 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s195  (
	.I0(\top/processor/sha_core/n327_169 ),
	.I1(\top/processor/sha_core/n327_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_199 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s196  (
	.I0(\top/processor/sha_core/n327_173 ),
	.I1(\top/processor/sha_core/n327_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_201 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s197  (
	.I0(\top/processor/sha_core/n327_177 ),
	.I1(\top/processor/sha_core/n327_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_203 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s198  (
	.I0(\top/processor/sha_core/n327_181 ),
	.I1(\top/processor/sha_core/n327_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_205 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s199  (
	.I0(\top/processor/sha_core/n327_185 ),
	.I1(\top/processor/sha_core/n327_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_207 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s200  (
	.I0(\top/processor/sha_core/n327_189 ),
	.I1(\top/processor/sha_core/n327_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_209 )
);
MUX2_LUT6 \top/processor/sha_core/n327_s201  (
	.I0(\top/processor/sha_core/n327_193 ),
	.I1(\top/processor/sha_core/n327_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n327_211 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s194  (
	.I0(\top/processor/sha_core/n328_165 ),
	.I1(\top/processor/sha_core/n328_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_197 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s195  (
	.I0(\top/processor/sha_core/n328_169 ),
	.I1(\top/processor/sha_core/n328_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_199 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s196  (
	.I0(\top/processor/sha_core/n328_173 ),
	.I1(\top/processor/sha_core/n328_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_201 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s197  (
	.I0(\top/processor/sha_core/n328_177 ),
	.I1(\top/processor/sha_core/n328_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_203 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s198  (
	.I0(\top/processor/sha_core/n328_181 ),
	.I1(\top/processor/sha_core/n328_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_205 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s199  (
	.I0(\top/processor/sha_core/n328_185 ),
	.I1(\top/processor/sha_core/n328_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_207 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s200  (
	.I0(\top/processor/sha_core/n328_189 ),
	.I1(\top/processor/sha_core/n328_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_209 )
);
MUX2_LUT6 \top/processor/sha_core/n328_s201  (
	.I0(\top/processor/sha_core/n328_193 ),
	.I1(\top/processor/sha_core/n328_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n328_211 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s194  (
	.I0(\top/processor/sha_core/n329_165 ),
	.I1(\top/processor/sha_core/n329_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_197 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s195  (
	.I0(\top/processor/sha_core/n329_169 ),
	.I1(\top/processor/sha_core/n329_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_199 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s196  (
	.I0(\top/processor/sha_core/n329_173 ),
	.I1(\top/processor/sha_core/n329_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_201 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s197  (
	.I0(\top/processor/sha_core/n329_177 ),
	.I1(\top/processor/sha_core/n329_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_203 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s198  (
	.I0(\top/processor/sha_core/n329_181 ),
	.I1(\top/processor/sha_core/n329_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_205 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s199  (
	.I0(\top/processor/sha_core/n329_185 ),
	.I1(\top/processor/sha_core/n329_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_207 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s200  (
	.I0(\top/processor/sha_core/n329_189 ),
	.I1(\top/processor/sha_core/n329_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_209 )
);
MUX2_LUT6 \top/processor/sha_core/n329_s201  (
	.I0(\top/processor/sha_core/n329_193 ),
	.I1(\top/processor/sha_core/n329_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n329_211 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s194  (
	.I0(\top/processor/sha_core/n330_165 ),
	.I1(\top/processor/sha_core/n330_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_197 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s195  (
	.I0(\top/processor/sha_core/n330_169 ),
	.I1(\top/processor/sha_core/n330_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_199 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s196  (
	.I0(\top/processor/sha_core/n330_173 ),
	.I1(\top/processor/sha_core/n330_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_201 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s197  (
	.I0(\top/processor/sha_core/n330_177 ),
	.I1(\top/processor/sha_core/n330_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_203 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s198  (
	.I0(\top/processor/sha_core/n330_181 ),
	.I1(\top/processor/sha_core/n330_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_205 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s199  (
	.I0(\top/processor/sha_core/n330_185 ),
	.I1(\top/processor/sha_core/n330_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_207 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s200  (
	.I0(\top/processor/sha_core/n330_189 ),
	.I1(\top/processor/sha_core/n330_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_209 )
);
MUX2_LUT6 \top/processor/sha_core/n330_s201  (
	.I0(\top/processor/sha_core/n330_193 ),
	.I1(\top/processor/sha_core/n330_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n330_211 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s194  (
	.I0(\top/processor/sha_core/n331_165 ),
	.I1(\top/processor/sha_core/n331_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_197 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s195  (
	.I0(\top/processor/sha_core/n331_169 ),
	.I1(\top/processor/sha_core/n331_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_199 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s196  (
	.I0(\top/processor/sha_core/n331_173 ),
	.I1(\top/processor/sha_core/n331_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_201 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s197  (
	.I0(\top/processor/sha_core/n331_177 ),
	.I1(\top/processor/sha_core/n331_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_203 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s198  (
	.I0(\top/processor/sha_core/n331_181 ),
	.I1(\top/processor/sha_core/n331_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_205 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s199  (
	.I0(\top/processor/sha_core/n331_185 ),
	.I1(\top/processor/sha_core/n331_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_207 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s200  (
	.I0(\top/processor/sha_core/n331_189 ),
	.I1(\top/processor/sha_core/n331_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_209 )
);
MUX2_LUT6 \top/processor/sha_core/n331_s201  (
	.I0(\top/processor/sha_core/n331_193 ),
	.I1(\top/processor/sha_core/n331_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n331_211 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s194  (
	.I0(\top/processor/sha_core/n332_165 ),
	.I1(\top/processor/sha_core/n332_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_197 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s195  (
	.I0(\top/processor/sha_core/n332_169 ),
	.I1(\top/processor/sha_core/n332_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_199 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s196  (
	.I0(\top/processor/sha_core/n332_173 ),
	.I1(\top/processor/sha_core/n332_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_201 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s197  (
	.I0(\top/processor/sha_core/n332_177 ),
	.I1(\top/processor/sha_core/n332_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_203 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s198  (
	.I0(\top/processor/sha_core/n332_181 ),
	.I1(\top/processor/sha_core/n332_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_205 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s199  (
	.I0(\top/processor/sha_core/n332_185 ),
	.I1(\top/processor/sha_core/n332_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_207 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s200  (
	.I0(\top/processor/sha_core/n332_189 ),
	.I1(\top/processor/sha_core/n332_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_209 )
);
MUX2_LUT6 \top/processor/sha_core/n332_s201  (
	.I0(\top/processor/sha_core/n332_193 ),
	.I1(\top/processor/sha_core/n332_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n332_211 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s194  (
	.I0(\top/processor/sha_core/n333_165 ),
	.I1(\top/processor/sha_core/n333_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_197 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s195  (
	.I0(\top/processor/sha_core/n333_169 ),
	.I1(\top/processor/sha_core/n333_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_199 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s196  (
	.I0(\top/processor/sha_core/n333_173 ),
	.I1(\top/processor/sha_core/n333_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_201 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s197  (
	.I0(\top/processor/sha_core/n333_177 ),
	.I1(\top/processor/sha_core/n333_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_203 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s198  (
	.I0(\top/processor/sha_core/n333_181 ),
	.I1(\top/processor/sha_core/n333_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_205 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s199  (
	.I0(\top/processor/sha_core/n333_185 ),
	.I1(\top/processor/sha_core/n333_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_207 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s200  (
	.I0(\top/processor/sha_core/n333_189 ),
	.I1(\top/processor/sha_core/n333_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_209 )
);
MUX2_LUT6 \top/processor/sha_core/n333_s201  (
	.I0(\top/processor/sha_core/n333_193 ),
	.I1(\top/processor/sha_core/n333_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n333_211 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s194  (
	.I0(\top/processor/sha_core/n334_165 ),
	.I1(\top/processor/sha_core/n334_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_197 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s195  (
	.I0(\top/processor/sha_core/n334_169 ),
	.I1(\top/processor/sha_core/n334_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_199 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s196  (
	.I0(\top/processor/sha_core/n334_173 ),
	.I1(\top/processor/sha_core/n334_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_201 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s197  (
	.I0(\top/processor/sha_core/n334_177 ),
	.I1(\top/processor/sha_core/n334_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_203 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s198  (
	.I0(\top/processor/sha_core/n334_181 ),
	.I1(\top/processor/sha_core/n334_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_205 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s199  (
	.I0(\top/processor/sha_core/n334_185 ),
	.I1(\top/processor/sha_core/n334_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_207 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s200  (
	.I0(\top/processor/sha_core/n334_189 ),
	.I1(\top/processor/sha_core/n334_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_209 )
);
MUX2_LUT6 \top/processor/sha_core/n334_s201  (
	.I0(\top/processor/sha_core/n334_193 ),
	.I1(\top/processor/sha_core/n334_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n334_211 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s194  (
	.I0(\top/processor/sha_core/n335_165 ),
	.I1(\top/processor/sha_core/n335_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_197 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s195  (
	.I0(\top/processor/sha_core/n335_169 ),
	.I1(\top/processor/sha_core/n335_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_199 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s196  (
	.I0(\top/processor/sha_core/n335_173 ),
	.I1(\top/processor/sha_core/n335_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_201 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s197  (
	.I0(\top/processor/sha_core/n335_177 ),
	.I1(\top/processor/sha_core/n335_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_203 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s198  (
	.I0(\top/processor/sha_core/n335_181 ),
	.I1(\top/processor/sha_core/n335_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_205 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s199  (
	.I0(\top/processor/sha_core/n335_185 ),
	.I1(\top/processor/sha_core/n335_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_207 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s200  (
	.I0(\top/processor/sha_core/n335_189 ),
	.I1(\top/processor/sha_core/n335_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_209 )
);
MUX2_LUT6 \top/processor/sha_core/n335_s201  (
	.I0(\top/processor/sha_core/n335_193 ),
	.I1(\top/processor/sha_core/n335_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n335_211 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s194  (
	.I0(\top/processor/sha_core/n336_165 ),
	.I1(\top/processor/sha_core/n336_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_197 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s195  (
	.I0(\top/processor/sha_core/n336_169 ),
	.I1(\top/processor/sha_core/n336_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_199 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s196  (
	.I0(\top/processor/sha_core/n336_173 ),
	.I1(\top/processor/sha_core/n336_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_201 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s197  (
	.I0(\top/processor/sha_core/n336_177 ),
	.I1(\top/processor/sha_core/n336_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_203 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s198  (
	.I0(\top/processor/sha_core/n336_181 ),
	.I1(\top/processor/sha_core/n336_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_205 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s199  (
	.I0(\top/processor/sha_core/n336_185 ),
	.I1(\top/processor/sha_core/n336_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_207 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s200  (
	.I0(\top/processor/sha_core/n336_189 ),
	.I1(\top/processor/sha_core/n336_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_209 )
);
MUX2_LUT6 \top/processor/sha_core/n336_s201  (
	.I0(\top/processor/sha_core/n336_193 ),
	.I1(\top/processor/sha_core/n336_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n336_211 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s194  (
	.I0(\top/processor/sha_core/n337_165 ),
	.I1(\top/processor/sha_core/n337_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_197 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s195  (
	.I0(\top/processor/sha_core/n337_169 ),
	.I1(\top/processor/sha_core/n337_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_199 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s196  (
	.I0(\top/processor/sha_core/n337_173 ),
	.I1(\top/processor/sha_core/n337_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_201 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s197  (
	.I0(\top/processor/sha_core/n337_177 ),
	.I1(\top/processor/sha_core/n337_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_203 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s198  (
	.I0(\top/processor/sha_core/n337_181 ),
	.I1(\top/processor/sha_core/n337_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_205 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s199  (
	.I0(\top/processor/sha_core/n337_185 ),
	.I1(\top/processor/sha_core/n337_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_207 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s200  (
	.I0(\top/processor/sha_core/n337_189 ),
	.I1(\top/processor/sha_core/n337_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_209 )
);
MUX2_LUT6 \top/processor/sha_core/n337_s201  (
	.I0(\top/processor/sha_core/n337_193 ),
	.I1(\top/processor/sha_core/n337_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n337_211 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s194  (
	.I0(\top/processor/sha_core/n338_165 ),
	.I1(\top/processor/sha_core/n338_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_197 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s195  (
	.I0(\top/processor/sha_core/n338_169 ),
	.I1(\top/processor/sha_core/n338_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_199 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s196  (
	.I0(\top/processor/sha_core/n338_173 ),
	.I1(\top/processor/sha_core/n338_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_201 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s197  (
	.I0(\top/processor/sha_core/n338_177 ),
	.I1(\top/processor/sha_core/n338_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_203 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s198  (
	.I0(\top/processor/sha_core/n338_181 ),
	.I1(\top/processor/sha_core/n338_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_205 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s199  (
	.I0(\top/processor/sha_core/n338_185 ),
	.I1(\top/processor/sha_core/n338_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_207 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s200  (
	.I0(\top/processor/sha_core/n338_189 ),
	.I1(\top/processor/sha_core/n338_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_209 )
);
MUX2_LUT6 \top/processor/sha_core/n338_s201  (
	.I0(\top/processor/sha_core/n338_193 ),
	.I1(\top/processor/sha_core/n338_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n338_211 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s194  (
	.I0(\top/processor/sha_core/n339_165 ),
	.I1(\top/processor/sha_core/n339_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_197 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s195  (
	.I0(\top/processor/sha_core/n339_169 ),
	.I1(\top/processor/sha_core/n339_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_199 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s196  (
	.I0(\top/processor/sha_core/n339_173 ),
	.I1(\top/processor/sha_core/n339_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_201 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s197  (
	.I0(\top/processor/sha_core/n339_177 ),
	.I1(\top/processor/sha_core/n339_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_203 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s198  (
	.I0(\top/processor/sha_core/n339_181 ),
	.I1(\top/processor/sha_core/n339_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_205 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s199  (
	.I0(\top/processor/sha_core/n339_185 ),
	.I1(\top/processor/sha_core/n339_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_207 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s200  (
	.I0(\top/processor/sha_core/n339_189 ),
	.I1(\top/processor/sha_core/n339_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_209 )
);
MUX2_LUT6 \top/processor/sha_core/n339_s201  (
	.I0(\top/processor/sha_core/n339_193 ),
	.I1(\top/processor/sha_core/n339_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n339_211 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s194  (
	.I0(\top/processor/sha_core/n340_165 ),
	.I1(\top/processor/sha_core/n340_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_197 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s195  (
	.I0(\top/processor/sha_core/n340_169 ),
	.I1(\top/processor/sha_core/n340_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_199 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s196  (
	.I0(\top/processor/sha_core/n340_173 ),
	.I1(\top/processor/sha_core/n340_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_201 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s197  (
	.I0(\top/processor/sha_core/n340_177 ),
	.I1(\top/processor/sha_core/n340_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_203 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s198  (
	.I0(\top/processor/sha_core/n340_181 ),
	.I1(\top/processor/sha_core/n340_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_205 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s199  (
	.I0(\top/processor/sha_core/n340_185 ),
	.I1(\top/processor/sha_core/n340_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_207 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s200  (
	.I0(\top/processor/sha_core/n340_189 ),
	.I1(\top/processor/sha_core/n340_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_209 )
);
MUX2_LUT6 \top/processor/sha_core/n340_s201  (
	.I0(\top/processor/sha_core/n340_193 ),
	.I1(\top/processor/sha_core/n340_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n340_211 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s194  (
	.I0(\top/processor/sha_core/n341_165 ),
	.I1(\top/processor/sha_core/n341_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_197 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s195  (
	.I0(\top/processor/sha_core/n341_169 ),
	.I1(\top/processor/sha_core/n341_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_199 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s196  (
	.I0(\top/processor/sha_core/n341_173 ),
	.I1(\top/processor/sha_core/n341_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_201 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s197  (
	.I0(\top/processor/sha_core/n341_177 ),
	.I1(\top/processor/sha_core/n341_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_203 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s198  (
	.I0(\top/processor/sha_core/n341_181 ),
	.I1(\top/processor/sha_core/n341_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_205 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s199  (
	.I0(\top/processor/sha_core/n341_185 ),
	.I1(\top/processor/sha_core/n341_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_207 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s200  (
	.I0(\top/processor/sha_core/n341_189 ),
	.I1(\top/processor/sha_core/n341_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_209 )
);
MUX2_LUT6 \top/processor/sha_core/n341_s201  (
	.I0(\top/processor/sha_core/n341_193 ),
	.I1(\top/processor/sha_core/n341_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n341_211 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s194  (
	.I0(\top/processor/sha_core/n342_165 ),
	.I1(\top/processor/sha_core/n342_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_197 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s195  (
	.I0(\top/processor/sha_core/n342_169 ),
	.I1(\top/processor/sha_core/n342_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_199 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s196  (
	.I0(\top/processor/sha_core/n342_173 ),
	.I1(\top/processor/sha_core/n342_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_201 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s197  (
	.I0(\top/processor/sha_core/n342_177 ),
	.I1(\top/processor/sha_core/n342_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_203 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s198  (
	.I0(\top/processor/sha_core/n342_181 ),
	.I1(\top/processor/sha_core/n342_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_205 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s199  (
	.I0(\top/processor/sha_core/n342_185 ),
	.I1(\top/processor/sha_core/n342_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_207 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s200  (
	.I0(\top/processor/sha_core/n342_189 ),
	.I1(\top/processor/sha_core/n342_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_209 )
);
MUX2_LUT6 \top/processor/sha_core/n342_s201  (
	.I0(\top/processor/sha_core/n342_193 ),
	.I1(\top/processor/sha_core/n342_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n342_211 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s194  (
	.I0(\top/processor/sha_core/n343_165 ),
	.I1(\top/processor/sha_core/n343_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_197 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s195  (
	.I0(\top/processor/sha_core/n343_169 ),
	.I1(\top/processor/sha_core/n343_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_199 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s196  (
	.I0(\top/processor/sha_core/n343_173 ),
	.I1(\top/processor/sha_core/n343_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_201 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s197  (
	.I0(\top/processor/sha_core/n343_177 ),
	.I1(\top/processor/sha_core/n343_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_203 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s198  (
	.I0(\top/processor/sha_core/n343_181 ),
	.I1(\top/processor/sha_core/n343_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_205 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s199  (
	.I0(\top/processor/sha_core/n343_185 ),
	.I1(\top/processor/sha_core/n343_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_207 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s200  (
	.I0(\top/processor/sha_core/n343_189 ),
	.I1(\top/processor/sha_core/n343_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_209 )
);
MUX2_LUT6 \top/processor/sha_core/n343_s201  (
	.I0(\top/processor/sha_core/n343_193 ),
	.I1(\top/processor/sha_core/n343_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n343_211 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s194  (
	.I0(\top/processor/sha_core/n344_165 ),
	.I1(\top/processor/sha_core/n344_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_197 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s195  (
	.I0(\top/processor/sha_core/n344_169 ),
	.I1(\top/processor/sha_core/n344_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_199 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s196  (
	.I0(\top/processor/sha_core/n344_173 ),
	.I1(\top/processor/sha_core/n344_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_201 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s197  (
	.I0(\top/processor/sha_core/n344_177 ),
	.I1(\top/processor/sha_core/n344_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_203 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s198  (
	.I0(\top/processor/sha_core/n344_181 ),
	.I1(\top/processor/sha_core/n344_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_205 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s199  (
	.I0(\top/processor/sha_core/n344_185 ),
	.I1(\top/processor/sha_core/n344_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_207 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s200  (
	.I0(\top/processor/sha_core/n344_189 ),
	.I1(\top/processor/sha_core/n344_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_209 )
);
MUX2_LUT6 \top/processor/sha_core/n344_s201  (
	.I0(\top/processor/sha_core/n344_193 ),
	.I1(\top/processor/sha_core/n344_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n344_211 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s194  (
	.I0(\top/processor/sha_core/n345_165 ),
	.I1(\top/processor/sha_core/n345_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_197 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s195  (
	.I0(\top/processor/sha_core/n345_169 ),
	.I1(\top/processor/sha_core/n345_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_199 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s196  (
	.I0(\top/processor/sha_core/n345_173 ),
	.I1(\top/processor/sha_core/n345_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_201 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s197  (
	.I0(\top/processor/sha_core/n345_177 ),
	.I1(\top/processor/sha_core/n345_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_203 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s198  (
	.I0(\top/processor/sha_core/n345_181 ),
	.I1(\top/processor/sha_core/n345_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_205 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s199  (
	.I0(\top/processor/sha_core/n345_185 ),
	.I1(\top/processor/sha_core/n345_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_207 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s200  (
	.I0(\top/processor/sha_core/n345_189 ),
	.I1(\top/processor/sha_core/n345_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_209 )
);
MUX2_LUT6 \top/processor/sha_core/n345_s201  (
	.I0(\top/processor/sha_core/n345_193 ),
	.I1(\top/processor/sha_core/n345_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n345_211 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s194  (
	.I0(\top/processor/sha_core/n346_165 ),
	.I1(\top/processor/sha_core/n346_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_197 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s195  (
	.I0(\top/processor/sha_core/n346_169 ),
	.I1(\top/processor/sha_core/n346_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_199 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s196  (
	.I0(\top/processor/sha_core/n346_173 ),
	.I1(\top/processor/sha_core/n346_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_201 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s197  (
	.I0(\top/processor/sha_core/n346_177 ),
	.I1(\top/processor/sha_core/n346_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_203 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s198  (
	.I0(\top/processor/sha_core/n346_181 ),
	.I1(\top/processor/sha_core/n346_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_205 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s199  (
	.I0(\top/processor/sha_core/n346_185 ),
	.I1(\top/processor/sha_core/n346_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_207 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s200  (
	.I0(\top/processor/sha_core/n346_189 ),
	.I1(\top/processor/sha_core/n346_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_209 )
);
MUX2_LUT6 \top/processor/sha_core/n346_s201  (
	.I0(\top/processor/sha_core/n346_193 ),
	.I1(\top/processor/sha_core/n346_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n346_211 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s194  (
	.I0(\top/processor/sha_core/n347_165 ),
	.I1(\top/processor/sha_core/n347_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_197 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s195  (
	.I0(\top/processor/sha_core/n347_169 ),
	.I1(\top/processor/sha_core/n347_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_199 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s196  (
	.I0(\top/processor/sha_core/n347_173 ),
	.I1(\top/processor/sha_core/n347_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_201 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s197  (
	.I0(\top/processor/sha_core/n347_177 ),
	.I1(\top/processor/sha_core/n347_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_203 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s198  (
	.I0(\top/processor/sha_core/n347_181 ),
	.I1(\top/processor/sha_core/n347_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_205 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s199  (
	.I0(\top/processor/sha_core/n347_185 ),
	.I1(\top/processor/sha_core/n347_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_207 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s200  (
	.I0(\top/processor/sha_core/n347_189 ),
	.I1(\top/processor/sha_core/n347_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_209 )
);
MUX2_LUT6 \top/processor/sha_core/n347_s201  (
	.I0(\top/processor/sha_core/n347_193 ),
	.I1(\top/processor/sha_core/n347_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n347_211 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s194  (
	.I0(\top/processor/sha_core/n348_165 ),
	.I1(\top/processor/sha_core/n348_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_197 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s195  (
	.I0(\top/processor/sha_core/n348_169 ),
	.I1(\top/processor/sha_core/n348_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_199 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s196  (
	.I0(\top/processor/sha_core/n348_173 ),
	.I1(\top/processor/sha_core/n348_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_201 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s197  (
	.I0(\top/processor/sha_core/n348_177 ),
	.I1(\top/processor/sha_core/n348_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_203 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s198  (
	.I0(\top/processor/sha_core/n348_181 ),
	.I1(\top/processor/sha_core/n348_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_205 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s199  (
	.I0(\top/processor/sha_core/n348_185 ),
	.I1(\top/processor/sha_core/n348_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_207 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s200  (
	.I0(\top/processor/sha_core/n348_189 ),
	.I1(\top/processor/sha_core/n348_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_209 )
);
MUX2_LUT6 \top/processor/sha_core/n348_s201  (
	.I0(\top/processor/sha_core/n348_193 ),
	.I1(\top/processor/sha_core/n348_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n348_211 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s194  (
	.I0(\top/processor/sha_core/n349_165 ),
	.I1(\top/processor/sha_core/n349_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_197 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s195  (
	.I0(\top/processor/sha_core/n349_169 ),
	.I1(\top/processor/sha_core/n349_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_199 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s196  (
	.I0(\top/processor/sha_core/n349_173 ),
	.I1(\top/processor/sha_core/n349_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_201 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s197  (
	.I0(\top/processor/sha_core/n349_177 ),
	.I1(\top/processor/sha_core/n349_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_203 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s198  (
	.I0(\top/processor/sha_core/n349_181 ),
	.I1(\top/processor/sha_core/n349_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_205 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s199  (
	.I0(\top/processor/sha_core/n349_185 ),
	.I1(\top/processor/sha_core/n349_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_207 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s200  (
	.I0(\top/processor/sha_core/n349_189 ),
	.I1(\top/processor/sha_core/n349_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_209 )
);
MUX2_LUT6 \top/processor/sha_core/n349_s201  (
	.I0(\top/processor/sha_core/n349_193 ),
	.I1(\top/processor/sha_core/n349_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n349_211 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s194  (
	.I0(\top/processor/sha_core/n350_165 ),
	.I1(\top/processor/sha_core/n350_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_197 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s195  (
	.I0(\top/processor/sha_core/n350_169 ),
	.I1(\top/processor/sha_core/n350_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_199 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s196  (
	.I0(\top/processor/sha_core/n350_173 ),
	.I1(\top/processor/sha_core/n350_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_201 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s197  (
	.I0(\top/processor/sha_core/n350_177 ),
	.I1(\top/processor/sha_core/n350_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_203 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s198  (
	.I0(\top/processor/sha_core/n350_181 ),
	.I1(\top/processor/sha_core/n350_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_205 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s199  (
	.I0(\top/processor/sha_core/n350_185 ),
	.I1(\top/processor/sha_core/n350_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_207 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s200  (
	.I0(\top/processor/sha_core/n350_189 ),
	.I1(\top/processor/sha_core/n350_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_209 )
);
MUX2_LUT6 \top/processor/sha_core/n350_s201  (
	.I0(\top/processor/sha_core/n350_193 ),
	.I1(\top/processor/sha_core/n350_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n350_211 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s194  (
	.I0(\top/processor/sha_core/n351_165 ),
	.I1(\top/processor/sha_core/n351_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_197 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s195  (
	.I0(\top/processor/sha_core/n351_169 ),
	.I1(\top/processor/sha_core/n351_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_199 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s196  (
	.I0(\top/processor/sha_core/n351_173 ),
	.I1(\top/processor/sha_core/n351_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_201 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s197  (
	.I0(\top/processor/sha_core/n351_177 ),
	.I1(\top/processor/sha_core/n351_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_203 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s198  (
	.I0(\top/processor/sha_core/n351_181 ),
	.I1(\top/processor/sha_core/n351_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_205 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s199  (
	.I0(\top/processor/sha_core/n351_185 ),
	.I1(\top/processor/sha_core/n351_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_207 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s200  (
	.I0(\top/processor/sha_core/n351_189 ),
	.I1(\top/processor/sha_core/n351_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_209 )
);
MUX2_LUT6 \top/processor/sha_core/n351_s201  (
	.I0(\top/processor/sha_core/n351_193 ),
	.I1(\top/processor/sha_core/n351_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n351_211 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s194  (
	.I0(\top/processor/sha_core/n352_165 ),
	.I1(\top/processor/sha_core/n352_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_197 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s195  (
	.I0(\top/processor/sha_core/n352_169 ),
	.I1(\top/processor/sha_core/n352_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_199 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s196  (
	.I0(\top/processor/sha_core/n352_173 ),
	.I1(\top/processor/sha_core/n352_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_201 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s197  (
	.I0(\top/processor/sha_core/n352_177 ),
	.I1(\top/processor/sha_core/n352_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_203 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s198  (
	.I0(\top/processor/sha_core/n352_181 ),
	.I1(\top/processor/sha_core/n352_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_205 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s199  (
	.I0(\top/processor/sha_core/n352_185 ),
	.I1(\top/processor/sha_core/n352_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_207 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s200  (
	.I0(\top/processor/sha_core/n352_189 ),
	.I1(\top/processor/sha_core/n352_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_209 )
);
MUX2_LUT6 \top/processor/sha_core/n352_s201  (
	.I0(\top/processor/sha_core/n352_193 ),
	.I1(\top/processor/sha_core/n352_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n352_211 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s194  (
	.I0(\top/processor/sha_core/n353_165 ),
	.I1(\top/processor/sha_core/n353_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_197 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s195  (
	.I0(\top/processor/sha_core/n353_169 ),
	.I1(\top/processor/sha_core/n353_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_199 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s196  (
	.I0(\top/processor/sha_core/n353_173 ),
	.I1(\top/processor/sha_core/n353_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_201 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s197  (
	.I0(\top/processor/sha_core/n353_177 ),
	.I1(\top/processor/sha_core/n353_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_203 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s198  (
	.I0(\top/processor/sha_core/n353_181 ),
	.I1(\top/processor/sha_core/n353_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_205 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s199  (
	.I0(\top/processor/sha_core/n353_185 ),
	.I1(\top/processor/sha_core/n353_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_207 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s200  (
	.I0(\top/processor/sha_core/n353_189 ),
	.I1(\top/processor/sha_core/n353_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_209 )
);
MUX2_LUT6 \top/processor/sha_core/n353_s201  (
	.I0(\top/processor/sha_core/n353_193 ),
	.I1(\top/processor/sha_core/n353_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n353_211 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s194  (
	.I0(\top/processor/sha_core/n354_165 ),
	.I1(\top/processor/sha_core/n354_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_197 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s195  (
	.I0(\top/processor/sha_core/n354_169 ),
	.I1(\top/processor/sha_core/n354_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_199 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s196  (
	.I0(\top/processor/sha_core/n354_173 ),
	.I1(\top/processor/sha_core/n354_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_201 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s197  (
	.I0(\top/processor/sha_core/n354_177 ),
	.I1(\top/processor/sha_core/n354_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_203 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s198  (
	.I0(\top/processor/sha_core/n354_181 ),
	.I1(\top/processor/sha_core/n354_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_205 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s199  (
	.I0(\top/processor/sha_core/n354_185 ),
	.I1(\top/processor/sha_core/n354_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_207 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s200  (
	.I0(\top/processor/sha_core/n354_189 ),
	.I1(\top/processor/sha_core/n354_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_209 )
);
MUX2_LUT6 \top/processor/sha_core/n354_s201  (
	.I0(\top/processor/sha_core/n354_193 ),
	.I1(\top/processor/sha_core/n354_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n354_211 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s194  (
	.I0(\top/processor/sha_core/n355_165 ),
	.I1(\top/processor/sha_core/n355_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_197 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s195  (
	.I0(\top/processor/sha_core/n355_169 ),
	.I1(\top/processor/sha_core/n355_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_199 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s196  (
	.I0(\top/processor/sha_core/n355_173 ),
	.I1(\top/processor/sha_core/n355_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_201 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s197  (
	.I0(\top/processor/sha_core/n355_177 ),
	.I1(\top/processor/sha_core/n355_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_203 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s198  (
	.I0(\top/processor/sha_core/n355_181 ),
	.I1(\top/processor/sha_core/n355_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_205 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s199  (
	.I0(\top/processor/sha_core/n355_185 ),
	.I1(\top/processor/sha_core/n355_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_207 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s200  (
	.I0(\top/processor/sha_core/n355_189 ),
	.I1(\top/processor/sha_core/n355_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_209 )
);
MUX2_LUT6 \top/processor/sha_core/n355_s201  (
	.I0(\top/processor/sha_core/n355_193 ),
	.I1(\top/processor/sha_core/n355_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n355_211 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s194  (
	.I0(\top/processor/sha_core/n356_165 ),
	.I1(\top/processor/sha_core/n356_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_197 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s195  (
	.I0(\top/processor/sha_core/n356_169 ),
	.I1(\top/processor/sha_core/n356_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_199 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s196  (
	.I0(\top/processor/sha_core/n356_173 ),
	.I1(\top/processor/sha_core/n356_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_201 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s197  (
	.I0(\top/processor/sha_core/n356_177 ),
	.I1(\top/processor/sha_core/n356_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_203 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s198  (
	.I0(\top/processor/sha_core/n356_181 ),
	.I1(\top/processor/sha_core/n356_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_205 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s199  (
	.I0(\top/processor/sha_core/n356_185 ),
	.I1(\top/processor/sha_core/n356_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_207 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s200  (
	.I0(\top/processor/sha_core/n356_189 ),
	.I1(\top/processor/sha_core/n356_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_209 )
);
MUX2_LUT6 \top/processor/sha_core/n356_s201  (
	.I0(\top/processor/sha_core/n356_193 ),
	.I1(\top/processor/sha_core/n356_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n356_211 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s194  (
	.I0(\top/processor/sha_core/n357_165 ),
	.I1(\top/processor/sha_core/n357_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_197 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s195  (
	.I0(\top/processor/sha_core/n357_169 ),
	.I1(\top/processor/sha_core/n357_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_199 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s196  (
	.I0(\top/processor/sha_core/n357_173 ),
	.I1(\top/processor/sha_core/n357_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_201 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s197  (
	.I0(\top/processor/sha_core/n357_177 ),
	.I1(\top/processor/sha_core/n357_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_203 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s198  (
	.I0(\top/processor/sha_core/n357_181 ),
	.I1(\top/processor/sha_core/n357_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_205 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s199  (
	.I0(\top/processor/sha_core/n357_185 ),
	.I1(\top/processor/sha_core/n357_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_207 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s200  (
	.I0(\top/processor/sha_core/n357_189 ),
	.I1(\top/processor/sha_core/n357_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_209 )
);
MUX2_LUT6 \top/processor/sha_core/n357_s201  (
	.I0(\top/processor/sha_core/n357_193 ),
	.I1(\top/processor/sha_core/n357_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n357_211 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s194  (
	.I0(\top/processor/sha_core/n358_165 ),
	.I1(\top/processor/sha_core/n358_167 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_197 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s195  (
	.I0(\top/processor/sha_core/n358_169 ),
	.I1(\top/processor/sha_core/n358_171 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_199 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s196  (
	.I0(\top/processor/sha_core/n358_173 ),
	.I1(\top/processor/sha_core/n358_175 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_201 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s197  (
	.I0(\top/processor/sha_core/n358_177 ),
	.I1(\top/processor/sha_core/n358_179 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_203 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s198  (
	.I0(\top/processor/sha_core/n358_181 ),
	.I1(\top/processor/sha_core/n358_183 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_205 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s199  (
	.I0(\top/processor/sha_core/n358_185 ),
	.I1(\top/processor/sha_core/n358_187 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_207 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s200  (
	.I0(\top/processor/sha_core/n358_189 ),
	.I1(\top/processor/sha_core/n358_191 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_209 )
);
MUX2_LUT6 \top/processor/sha_core/n358_s201  (
	.I0(\top/processor/sha_core/n358_193 ),
	.I1(\top/processor/sha_core/n358_195 ),
	.S0(\top/processor/sha_core/t [2]),
	.O(\top/processor/sha_core/n358_211 )
);
MUX2_LUT6 \top/processor/sha_core/n3488_s174  (
	.I0(\top/processor/sha_core/n3488_181 ),
	.I1(\top/processor/sha_core/n3488_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3488_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3488_s175  (
	.I0(\top/processor/sha_core/n3488_185 ),
	.I1(\top/processor/sha_core/n3488_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3488_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3489_s174  (
	.I0(\top/processor/sha_core/n3489_181 ),
	.I1(\top/processor/sha_core/n3489_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3489_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3489_s175  (
	.I0(\top/processor/sha_core/n3489_185 ),
	.I1(\top/processor/sha_core/n3489_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3489_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3490_s174  (
	.I0(\top/processor/sha_core/n3490_181 ),
	.I1(\top/processor/sha_core/n3490_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3490_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3490_s175  (
	.I0(\top/processor/sha_core/n3490_185 ),
	.I1(\top/processor/sha_core/n3490_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3490_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3491_s174  (
	.I0(\top/processor/sha_core/n3491_181 ),
	.I1(\top/processor/sha_core/n3491_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3491_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3491_s175  (
	.I0(\top/processor/sha_core/n3491_185 ),
	.I1(\top/processor/sha_core/n3491_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3491_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3492_s174  (
	.I0(\top/processor/sha_core/n3492_181 ),
	.I1(\top/processor/sha_core/n3492_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3492_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3492_s175  (
	.I0(\top/processor/sha_core/n3492_185 ),
	.I1(\top/processor/sha_core/n3492_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3492_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3493_s174  (
	.I0(\top/processor/sha_core/n3493_181 ),
	.I1(\top/processor/sha_core/n3493_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3493_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3493_s175  (
	.I0(\top/processor/sha_core/n3493_185 ),
	.I1(\top/processor/sha_core/n3493_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3493_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3494_s174  (
	.I0(\top/processor/sha_core/n3494_182 ),
	.I1(\top/processor/sha_core/n3494_184 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3494_190 )
);
MUX2_LUT6 \top/processor/sha_core/n3494_s175  (
	.I0(\top/processor/sha_core/n3494_186 ),
	.I1(\top/processor/sha_core/n3494_188 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3494_192 )
);
MUX2_LUT6 \top/processor/sha_core/n3495_s174  (
	.I0(\top/processor/sha_core/n3495_181 ),
	.I1(\top/processor/sha_core/n3495_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3495_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3495_s175  (
	.I0(\top/processor/sha_core/n3495_185 ),
	.I1(\top/processor/sha_core/n3495_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3495_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3496_s174  (
	.I0(\top/processor/sha_core/n3496_181 ),
	.I1(\top/processor/sha_core/n3496_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3496_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3496_s175  (
	.I0(\top/processor/sha_core/n3496_185 ),
	.I1(\top/processor/sha_core/n3496_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3496_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3497_s174  (
	.I0(\top/processor/sha_core/n3497_181 ),
	.I1(\top/processor/sha_core/n3497_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3497_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3497_s175  (
	.I0(\top/processor/sha_core/n3497_185 ),
	.I1(\top/processor/sha_core/n3497_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3497_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3498_s174  (
	.I0(\top/processor/sha_core/n3498_181 ),
	.I1(\top/processor/sha_core/n3498_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3498_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3498_s175  (
	.I0(\top/processor/sha_core/n3498_185 ),
	.I1(\top/processor/sha_core/n3498_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3498_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3499_s174  (
	.I0(\top/processor/sha_core/n3499_181 ),
	.I1(\top/processor/sha_core/n3499_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3499_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3499_s175  (
	.I0(\top/processor/sha_core/n3499_185 ),
	.I1(\top/processor/sha_core/n3499_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3499_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3500_s174  (
	.I0(\top/processor/sha_core/n3500_181 ),
	.I1(\top/processor/sha_core/n3500_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3500_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3500_s175  (
	.I0(\top/processor/sha_core/n3500_185 ),
	.I1(\top/processor/sha_core/n3500_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3500_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3501_s174  (
	.I0(\top/processor/sha_core/n3501_181 ),
	.I1(\top/processor/sha_core/n3501_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3501_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3501_s175  (
	.I0(\top/processor/sha_core/n3501_185 ),
	.I1(\top/processor/sha_core/n3501_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3501_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3502_s174  (
	.I0(\top/processor/sha_core/n3502_181 ),
	.I1(\top/processor/sha_core/n3502_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3502_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3502_s175  (
	.I0(\top/processor/sha_core/n3502_185 ),
	.I1(\top/processor/sha_core/n3502_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3502_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3503_s174  (
	.I0(\top/processor/sha_core/n3503_181 ),
	.I1(\top/processor/sha_core/n3503_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3503_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3503_s175  (
	.I0(\top/processor/sha_core/n3503_185 ),
	.I1(\top/processor/sha_core/n3503_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3503_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3504_s174  (
	.I0(\top/processor/sha_core/n3504_181 ),
	.I1(\top/processor/sha_core/n3504_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3504_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3504_s175  (
	.I0(\top/processor/sha_core/n3504_185 ),
	.I1(\top/processor/sha_core/n3504_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3504_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3505_s174  (
	.I0(\top/processor/sha_core/n3505_181 ),
	.I1(\top/processor/sha_core/n3505_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3505_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3505_s175  (
	.I0(\top/processor/sha_core/n3505_185 ),
	.I1(\top/processor/sha_core/n3505_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3505_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3506_s174  (
	.I0(\top/processor/sha_core/n3506_181 ),
	.I1(\top/processor/sha_core/n3506_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3506_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3506_s175  (
	.I0(\top/processor/sha_core/n3506_185 ),
	.I1(\top/processor/sha_core/n3506_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3506_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3507_s174  (
	.I0(\top/processor/sha_core/n3507_181 ),
	.I1(\top/processor/sha_core/n3507_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3507_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3507_s175  (
	.I0(\top/processor/sha_core/n3507_185 ),
	.I1(\top/processor/sha_core/n3507_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3507_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3508_s174  (
	.I0(\top/processor/sha_core/n3508_181 ),
	.I1(\top/processor/sha_core/n3508_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3508_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3508_s175  (
	.I0(\top/processor/sha_core/n3508_185 ),
	.I1(\top/processor/sha_core/n3508_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3508_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3509_s174  (
	.I0(\top/processor/sha_core/n3509_181 ),
	.I1(\top/processor/sha_core/n3509_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3509_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3509_s175  (
	.I0(\top/processor/sha_core/n3509_185 ),
	.I1(\top/processor/sha_core/n3509_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3509_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3510_s171  (
	.I0(\top/processor/sha_core/n3510_181 ),
	.I1(\top/processor/sha_core/n3510_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3510_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3510_s172  (
	.I0(\top/processor/sha_core/n3510_185 ),
	.I1(\top/processor/sha_core/n3510_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3510_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3511_s174  (
	.I0(\top/processor/sha_core/n3511_181 ),
	.I1(\top/processor/sha_core/n3511_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3511_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3511_s175  (
	.I0(\top/processor/sha_core/n3511_185 ),
	.I1(\top/processor/sha_core/n3511_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3511_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3512_s174  (
	.I0(\top/processor/sha_core/n3512_181 ),
	.I1(\top/processor/sha_core/n3512_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3512_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3512_s175  (
	.I0(\top/processor/sha_core/n3512_185 ),
	.I1(\top/processor/sha_core/n3512_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3512_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3513_s174  (
	.I0(\top/processor/sha_core/n3513_181 ),
	.I1(\top/processor/sha_core/n3513_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3513_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3513_s175  (
	.I0(\top/processor/sha_core/n3513_185 ),
	.I1(\top/processor/sha_core/n3513_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3513_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3514_s174  (
	.I0(\top/processor/sha_core/n3514_181 ),
	.I1(\top/processor/sha_core/n3514_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3514_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3514_s175  (
	.I0(\top/processor/sha_core/n3514_185 ),
	.I1(\top/processor/sha_core/n3514_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3514_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3515_s174  (
	.I0(\top/processor/sha_core/n3515_181 ),
	.I1(\top/processor/sha_core/n3515_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3515_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3515_s175  (
	.I0(\top/processor/sha_core/n3515_185 ),
	.I1(\top/processor/sha_core/n3515_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3515_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3516_s174  (
	.I0(\top/processor/sha_core/n3516_181 ),
	.I1(\top/processor/sha_core/n3516_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3516_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3516_s175  (
	.I0(\top/processor/sha_core/n3516_185 ),
	.I1(\top/processor/sha_core/n3516_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3516_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3517_s174  (
	.I0(\top/processor/sha_core/n3517_181 ),
	.I1(\top/processor/sha_core/n3517_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3517_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3517_s175  (
	.I0(\top/processor/sha_core/n3517_185 ),
	.I1(\top/processor/sha_core/n3517_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3517_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3518_s174  (
	.I0(\top/processor/sha_core/n3518_181 ),
	.I1(\top/processor/sha_core/n3518_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3518_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3518_s175  (
	.I0(\top/processor/sha_core/n3518_185 ),
	.I1(\top/processor/sha_core/n3518_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3518_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3519_s174  (
	.I0(\top/processor/sha_core/n3519_181 ),
	.I1(\top/processor/sha_core/n3519_183 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3519_189 )
);
MUX2_LUT6 \top/processor/sha_core/n3519_s175  (
	.I0(\top/processor/sha_core/n3519_185 ),
	.I1(\top/processor/sha_core/n3519_187 ),
	.S0(\top/processor/sha_core/n3460_11 ),
	.O(\top/processor/sha_core/n3519_191 )
);
MUX2_LUT6 \top/processor/sha_core/n3860_s126  (
	.I0(\top/processor/sha_core/n3860_135 ),
	.I1(\top/processor/sha_core/n3860_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3860_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3860_s127  (
	.I0(\top/processor/sha_core/n3860_139 ),
	.I1(\top/processor/sha_core/n3860_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3860_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3861_s126  (
	.I0(\top/processor/sha_core/n3861_135 ),
	.I1(\top/processor/sha_core/n3861_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3861_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3861_s127  (
	.I0(\top/processor/sha_core/n3861_139 ),
	.I1(\top/processor/sha_core/n3861_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3861_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3862_s126  (
	.I0(\top/processor/sha_core/n3862_135 ),
	.I1(\top/processor/sha_core/n3862_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3862_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3862_s127  (
	.I0(\top/processor/sha_core/n3862_139 ),
	.I1(\top/processor/sha_core/n3862_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3862_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3863_s126  (
	.I0(\top/processor/sha_core/n3863_135 ),
	.I1(\top/processor/sha_core/n3863_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3863_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3863_s127  (
	.I0(\top/processor/sha_core/n3863_139 ),
	.I1(\top/processor/sha_core/n3863_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3863_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3864_s126  (
	.I0(\top/processor/sha_core/n3864_135 ),
	.I1(\top/processor/sha_core/n3864_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3864_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3864_s127  (
	.I0(\top/processor/sha_core/n3864_139 ),
	.I1(\top/processor/sha_core/n3864_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3864_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3865_s126  (
	.I0(\top/processor/sha_core/n3865_135 ),
	.I1(\top/processor/sha_core/n3865_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3865_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3865_s127  (
	.I0(\top/processor/sha_core/n3865_139 ),
	.I1(\top/processor/sha_core/n3865_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3865_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3866_s126  (
	.I0(\top/processor/sha_core/n3866_135 ),
	.I1(\top/processor/sha_core/n3866_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3866_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3866_s127  (
	.I0(\top/processor/sha_core/n3866_139 ),
	.I1(\top/processor/sha_core/n3866_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3866_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3867_s126  (
	.I0(\top/processor/sha_core/n3867_135 ),
	.I1(\top/processor/sha_core/n3867_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3867_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3867_s127  (
	.I0(\top/processor/sha_core/n3867_139 ),
	.I1(\top/processor/sha_core/n3867_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3867_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3868_s126  (
	.I0(\top/processor/sha_core/n3868_135 ),
	.I1(\top/processor/sha_core/n3868_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3868_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3868_s127  (
	.I0(\top/processor/sha_core/n3868_139 ),
	.I1(\top/processor/sha_core/n3868_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3868_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3869_s126  (
	.I0(\top/processor/sha_core/n3869_135 ),
	.I1(\top/processor/sha_core/n3869_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3869_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3869_s127  (
	.I0(\top/processor/sha_core/n3869_139 ),
	.I1(\top/processor/sha_core/n3869_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3869_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3870_s126  (
	.I0(\top/processor/sha_core/n3870_135 ),
	.I1(\top/processor/sha_core/n3870_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3870_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3870_s127  (
	.I0(\top/processor/sha_core/n3870_139 ),
	.I1(\top/processor/sha_core/n3870_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3870_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3871_s126  (
	.I0(\top/processor/sha_core/n3871_135 ),
	.I1(\top/processor/sha_core/n3871_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3871_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3871_s127  (
	.I0(\top/processor/sha_core/n3871_139 ),
	.I1(\top/processor/sha_core/n3871_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3871_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3872_s126  (
	.I0(\top/processor/sha_core/n3872_135 ),
	.I1(\top/processor/sha_core/n3872_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3872_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3872_s127  (
	.I0(\top/processor/sha_core/n3872_139 ),
	.I1(\top/processor/sha_core/n3872_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3872_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3873_s126  (
	.I0(\top/processor/sha_core/n3873_135 ),
	.I1(\top/processor/sha_core/n3873_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3873_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3873_s127  (
	.I0(\top/processor/sha_core/n3873_139 ),
	.I1(\top/processor/sha_core/n3873_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3873_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3874_s126  (
	.I0(\top/processor/sha_core/n3874_135 ),
	.I1(\top/processor/sha_core/n3874_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3874_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3874_s127  (
	.I0(\top/processor/sha_core/n3874_139 ),
	.I1(\top/processor/sha_core/n3874_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3874_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3875_s126  (
	.I0(\top/processor/sha_core/n3875_135 ),
	.I1(\top/processor/sha_core/n3875_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3875_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3875_s127  (
	.I0(\top/processor/sha_core/n3875_139 ),
	.I1(\top/processor/sha_core/n3875_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3875_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3876_s126  (
	.I0(\top/processor/sha_core/n3876_135 ),
	.I1(\top/processor/sha_core/n3876_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3876_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3876_s127  (
	.I0(\top/processor/sha_core/n3876_139 ),
	.I1(\top/processor/sha_core/n3876_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3876_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3877_s126  (
	.I0(\top/processor/sha_core/n3877_135 ),
	.I1(\top/processor/sha_core/n3877_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3877_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3877_s127  (
	.I0(\top/processor/sha_core/n3877_139 ),
	.I1(\top/processor/sha_core/n3877_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3877_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3878_s126  (
	.I0(\top/processor/sha_core/n3878_135 ),
	.I1(\top/processor/sha_core/n3878_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3878_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3878_s127  (
	.I0(\top/processor/sha_core/n3878_139 ),
	.I1(\top/processor/sha_core/n3878_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3878_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3879_s126  (
	.I0(\top/processor/sha_core/n3879_135 ),
	.I1(\top/processor/sha_core/n3879_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3879_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3879_s127  (
	.I0(\top/processor/sha_core/n3879_139 ),
	.I1(\top/processor/sha_core/n3879_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3879_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3880_s126  (
	.I0(\top/processor/sha_core/n3880_135 ),
	.I1(\top/processor/sha_core/n3880_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3880_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3880_s127  (
	.I0(\top/processor/sha_core/n3880_139 ),
	.I1(\top/processor/sha_core/n3880_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3880_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3881_s126  (
	.I0(\top/processor/sha_core/n3881_135 ),
	.I1(\top/processor/sha_core/n3881_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3881_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3881_s127  (
	.I0(\top/processor/sha_core/n3881_139 ),
	.I1(\top/processor/sha_core/n3881_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3881_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3882_s126  (
	.I0(\top/processor/sha_core/n3882_135 ),
	.I1(\top/processor/sha_core/n3882_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3882_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3882_s127  (
	.I0(\top/processor/sha_core/n3882_139 ),
	.I1(\top/processor/sha_core/n3882_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3882_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3883_s126  (
	.I0(\top/processor/sha_core/n3883_135 ),
	.I1(\top/processor/sha_core/n3883_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3883_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3883_s127  (
	.I0(\top/processor/sha_core/n3883_139 ),
	.I1(\top/processor/sha_core/n3883_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3883_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3884_s126  (
	.I0(\top/processor/sha_core/n3884_135 ),
	.I1(\top/processor/sha_core/n3884_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3884_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3884_s127  (
	.I0(\top/processor/sha_core/n3884_139 ),
	.I1(\top/processor/sha_core/n3884_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3884_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3885_s126  (
	.I0(\top/processor/sha_core/n3885_135 ),
	.I1(\top/processor/sha_core/n3885_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3885_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3885_s127  (
	.I0(\top/processor/sha_core/n3885_139 ),
	.I1(\top/processor/sha_core/n3885_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3885_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3886_s126  (
	.I0(\top/processor/sha_core/n3886_135 ),
	.I1(\top/processor/sha_core/n3886_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3886_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3886_s127  (
	.I0(\top/processor/sha_core/n3886_139 ),
	.I1(\top/processor/sha_core/n3886_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3886_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3887_s126  (
	.I0(\top/processor/sha_core/n3887_135 ),
	.I1(\top/processor/sha_core/n3887_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3887_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3887_s127  (
	.I0(\top/processor/sha_core/n3887_139 ),
	.I1(\top/processor/sha_core/n3887_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3887_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3888_s126  (
	.I0(\top/processor/sha_core/n3888_135 ),
	.I1(\top/processor/sha_core/n3888_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3888_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3888_s127  (
	.I0(\top/processor/sha_core/n3888_139 ),
	.I1(\top/processor/sha_core/n3888_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3888_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3889_s126  (
	.I0(\top/processor/sha_core/n3889_135 ),
	.I1(\top/processor/sha_core/n3889_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3889_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3889_s127  (
	.I0(\top/processor/sha_core/n3889_139 ),
	.I1(\top/processor/sha_core/n3889_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3889_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3890_s126  (
	.I0(\top/processor/sha_core/n3890_135 ),
	.I1(\top/processor/sha_core/n3890_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3890_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3890_s127  (
	.I0(\top/processor/sha_core/n3890_139 ),
	.I1(\top/processor/sha_core/n3890_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3890_143 )
);
MUX2_LUT6 \top/processor/sha_core/n3891_s126  (
	.I0(\top/processor/sha_core/n3891_135 ),
	.I1(\top/processor/sha_core/n3891_133 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3891_141 )
);
MUX2_LUT6 \top/processor/sha_core/n3891_s127  (
	.I0(\top/processor/sha_core/n3891_139 ),
	.I1(\top/processor/sha_core/n3891_137 ),
	.S0(\top/processor/sha_core/msg_idx [4]),
	.O(\top/processor/sha_core/n3891_143 )
);
MUX2_LUT7 \top/processor/sha_core/n327_s190  (
	.I0(\top/processor/sha_core/n327_197 ),
	.I1(\top/processor/sha_core/n327_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n327_213 )
);
MUX2_LUT7 \top/processor/sha_core/n327_s191  (
	.I0(\top/processor/sha_core/n327_201 ),
	.I1(\top/processor/sha_core/n327_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n327_215 )
);
MUX2_LUT7 \top/processor/sha_core/n327_s192  (
	.I0(\top/processor/sha_core/n327_205 ),
	.I1(\top/processor/sha_core/n327_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n327_217 )
);
MUX2_LUT7 \top/processor/sha_core/n327_s193  (
	.I0(\top/processor/sha_core/n327_209 ),
	.I1(\top/processor/sha_core/n327_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n327_219 )
);
MUX2_LUT7 \top/processor/sha_core/n328_s190  (
	.I0(\top/processor/sha_core/n328_197 ),
	.I1(\top/processor/sha_core/n328_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n328_213 )
);
MUX2_LUT7 \top/processor/sha_core/n328_s191  (
	.I0(\top/processor/sha_core/n328_201 ),
	.I1(\top/processor/sha_core/n328_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n328_215 )
);
MUX2_LUT7 \top/processor/sha_core/n328_s192  (
	.I0(\top/processor/sha_core/n328_205 ),
	.I1(\top/processor/sha_core/n328_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n328_217 )
);
MUX2_LUT7 \top/processor/sha_core/n328_s193  (
	.I0(\top/processor/sha_core/n328_209 ),
	.I1(\top/processor/sha_core/n328_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n328_219 )
);
MUX2_LUT7 \top/processor/sha_core/n329_s190  (
	.I0(\top/processor/sha_core/n329_197 ),
	.I1(\top/processor/sha_core/n329_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n329_213 )
);
MUX2_LUT7 \top/processor/sha_core/n329_s191  (
	.I0(\top/processor/sha_core/n329_201 ),
	.I1(\top/processor/sha_core/n329_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n329_215 )
);
MUX2_LUT7 \top/processor/sha_core/n329_s192  (
	.I0(\top/processor/sha_core/n329_205 ),
	.I1(\top/processor/sha_core/n329_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n329_217 )
);
MUX2_LUT7 \top/processor/sha_core/n329_s193  (
	.I0(\top/processor/sha_core/n329_209 ),
	.I1(\top/processor/sha_core/n329_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n329_219 )
);
MUX2_LUT7 \top/processor/sha_core/n330_s190  (
	.I0(\top/processor/sha_core/n330_197 ),
	.I1(\top/processor/sha_core/n330_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n330_213 )
);
MUX2_LUT7 \top/processor/sha_core/n330_s191  (
	.I0(\top/processor/sha_core/n330_201 ),
	.I1(\top/processor/sha_core/n330_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n330_215 )
);
MUX2_LUT7 \top/processor/sha_core/n330_s192  (
	.I0(\top/processor/sha_core/n330_205 ),
	.I1(\top/processor/sha_core/n330_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n330_217 )
);
MUX2_LUT7 \top/processor/sha_core/n330_s193  (
	.I0(\top/processor/sha_core/n330_209 ),
	.I1(\top/processor/sha_core/n330_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n330_219 )
);
MUX2_LUT7 \top/processor/sha_core/n331_s190  (
	.I0(\top/processor/sha_core/n331_197 ),
	.I1(\top/processor/sha_core/n331_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n331_213 )
);
MUX2_LUT7 \top/processor/sha_core/n331_s191  (
	.I0(\top/processor/sha_core/n331_201 ),
	.I1(\top/processor/sha_core/n331_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n331_215 )
);
MUX2_LUT7 \top/processor/sha_core/n331_s192  (
	.I0(\top/processor/sha_core/n331_205 ),
	.I1(\top/processor/sha_core/n331_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n331_217 )
);
MUX2_LUT7 \top/processor/sha_core/n331_s193  (
	.I0(\top/processor/sha_core/n331_209 ),
	.I1(\top/processor/sha_core/n331_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n331_219 )
);
MUX2_LUT7 \top/processor/sha_core/n332_s190  (
	.I0(\top/processor/sha_core/n332_197 ),
	.I1(\top/processor/sha_core/n332_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n332_213 )
);
MUX2_LUT7 \top/processor/sha_core/n332_s191  (
	.I0(\top/processor/sha_core/n332_201 ),
	.I1(\top/processor/sha_core/n332_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n332_215 )
);
MUX2_LUT7 \top/processor/sha_core/n332_s192  (
	.I0(\top/processor/sha_core/n332_205 ),
	.I1(\top/processor/sha_core/n332_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n332_217 )
);
MUX2_LUT7 \top/processor/sha_core/n332_s193  (
	.I0(\top/processor/sha_core/n332_209 ),
	.I1(\top/processor/sha_core/n332_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n332_219 )
);
MUX2_LUT7 \top/processor/sha_core/n333_s190  (
	.I0(\top/processor/sha_core/n333_197 ),
	.I1(\top/processor/sha_core/n333_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n333_213 )
);
MUX2_LUT7 \top/processor/sha_core/n333_s191  (
	.I0(\top/processor/sha_core/n333_201 ),
	.I1(\top/processor/sha_core/n333_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n333_215 )
);
MUX2_LUT7 \top/processor/sha_core/n333_s192  (
	.I0(\top/processor/sha_core/n333_205 ),
	.I1(\top/processor/sha_core/n333_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n333_217 )
);
MUX2_LUT7 \top/processor/sha_core/n333_s193  (
	.I0(\top/processor/sha_core/n333_209 ),
	.I1(\top/processor/sha_core/n333_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n333_219 )
);
MUX2_LUT7 \top/processor/sha_core/n334_s190  (
	.I0(\top/processor/sha_core/n334_197 ),
	.I1(\top/processor/sha_core/n334_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n334_213 )
);
MUX2_LUT7 \top/processor/sha_core/n334_s191  (
	.I0(\top/processor/sha_core/n334_201 ),
	.I1(\top/processor/sha_core/n334_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n334_215 )
);
MUX2_LUT7 \top/processor/sha_core/n334_s192  (
	.I0(\top/processor/sha_core/n334_205 ),
	.I1(\top/processor/sha_core/n334_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n334_217 )
);
MUX2_LUT7 \top/processor/sha_core/n334_s193  (
	.I0(\top/processor/sha_core/n334_209 ),
	.I1(\top/processor/sha_core/n334_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n334_219 )
);
MUX2_LUT7 \top/processor/sha_core/n335_s190  (
	.I0(\top/processor/sha_core/n335_197 ),
	.I1(\top/processor/sha_core/n335_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n335_213 )
);
MUX2_LUT7 \top/processor/sha_core/n335_s191  (
	.I0(\top/processor/sha_core/n335_201 ),
	.I1(\top/processor/sha_core/n335_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n335_215 )
);
MUX2_LUT7 \top/processor/sha_core/n335_s192  (
	.I0(\top/processor/sha_core/n335_205 ),
	.I1(\top/processor/sha_core/n335_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n335_217 )
);
MUX2_LUT7 \top/processor/sha_core/n335_s193  (
	.I0(\top/processor/sha_core/n335_209 ),
	.I1(\top/processor/sha_core/n335_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n335_219 )
);
MUX2_LUT7 \top/processor/sha_core/n336_s190  (
	.I0(\top/processor/sha_core/n336_197 ),
	.I1(\top/processor/sha_core/n336_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n336_213 )
);
MUX2_LUT7 \top/processor/sha_core/n336_s191  (
	.I0(\top/processor/sha_core/n336_201 ),
	.I1(\top/processor/sha_core/n336_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n336_215 )
);
MUX2_LUT7 \top/processor/sha_core/n336_s192  (
	.I0(\top/processor/sha_core/n336_205 ),
	.I1(\top/processor/sha_core/n336_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n336_217 )
);
MUX2_LUT7 \top/processor/sha_core/n336_s193  (
	.I0(\top/processor/sha_core/n336_209 ),
	.I1(\top/processor/sha_core/n336_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n336_219 )
);
MUX2_LUT7 \top/processor/sha_core/n337_s190  (
	.I0(\top/processor/sha_core/n337_197 ),
	.I1(\top/processor/sha_core/n337_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n337_213 )
);
MUX2_LUT7 \top/processor/sha_core/n337_s191  (
	.I0(\top/processor/sha_core/n337_201 ),
	.I1(\top/processor/sha_core/n337_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n337_215 )
);
MUX2_LUT7 \top/processor/sha_core/n337_s192  (
	.I0(\top/processor/sha_core/n337_205 ),
	.I1(\top/processor/sha_core/n337_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n337_217 )
);
MUX2_LUT7 \top/processor/sha_core/n337_s193  (
	.I0(\top/processor/sha_core/n337_209 ),
	.I1(\top/processor/sha_core/n337_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n337_219 )
);
MUX2_LUT7 \top/processor/sha_core/n338_s190  (
	.I0(\top/processor/sha_core/n338_197 ),
	.I1(\top/processor/sha_core/n338_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n338_213 )
);
MUX2_LUT7 \top/processor/sha_core/n338_s191  (
	.I0(\top/processor/sha_core/n338_201 ),
	.I1(\top/processor/sha_core/n338_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n338_215 )
);
MUX2_LUT7 \top/processor/sha_core/n338_s192  (
	.I0(\top/processor/sha_core/n338_205 ),
	.I1(\top/processor/sha_core/n338_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n338_217 )
);
MUX2_LUT7 \top/processor/sha_core/n338_s193  (
	.I0(\top/processor/sha_core/n338_209 ),
	.I1(\top/processor/sha_core/n338_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n338_219 )
);
MUX2_LUT7 \top/processor/sha_core/n339_s190  (
	.I0(\top/processor/sha_core/n339_197 ),
	.I1(\top/processor/sha_core/n339_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n339_213 )
);
MUX2_LUT7 \top/processor/sha_core/n339_s191  (
	.I0(\top/processor/sha_core/n339_201 ),
	.I1(\top/processor/sha_core/n339_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n339_215 )
);
MUX2_LUT7 \top/processor/sha_core/n339_s192  (
	.I0(\top/processor/sha_core/n339_205 ),
	.I1(\top/processor/sha_core/n339_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n339_217 )
);
MUX2_LUT7 \top/processor/sha_core/n339_s193  (
	.I0(\top/processor/sha_core/n339_209 ),
	.I1(\top/processor/sha_core/n339_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n339_219 )
);
MUX2_LUT7 \top/processor/sha_core/n340_s190  (
	.I0(\top/processor/sha_core/n340_197 ),
	.I1(\top/processor/sha_core/n340_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n340_213 )
);
MUX2_LUT7 \top/processor/sha_core/n340_s191  (
	.I0(\top/processor/sha_core/n340_201 ),
	.I1(\top/processor/sha_core/n340_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n340_215 )
);
MUX2_LUT7 \top/processor/sha_core/n340_s192  (
	.I0(\top/processor/sha_core/n340_205 ),
	.I1(\top/processor/sha_core/n340_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n340_217 )
);
MUX2_LUT7 \top/processor/sha_core/n340_s193  (
	.I0(\top/processor/sha_core/n340_209 ),
	.I1(\top/processor/sha_core/n340_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n340_219 )
);
MUX2_LUT7 \top/processor/sha_core/n341_s190  (
	.I0(\top/processor/sha_core/n341_197 ),
	.I1(\top/processor/sha_core/n341_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n341_213 )
);
MUX2_LUT7 \top/processor/sha_core/n341_s191  (
	.I0(\top/processor/sha_core/n341_201 ),
	.I1(\top/processor/sha_core/n341_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n341_215 )
);
MUX2_LUT7 \top/processor/sha_core/n341_s192  (
	.I0(\top/processor/sha_core/n341_205 ),
	.I1(\top/processor/sha_core/n341_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n341_217 )
);
MUX2_LUT7 \top/processor/sha_core/n341_s193  (
	.I0(\top/processor/sha_core/n341_209 ),
	.I1(\top/processor/sha_core/n341_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n341_219 )
);
MUX2_LUT7 \top/processor/sha_core/n342_s190  (
	.I0(\top/processor/sha_core/n342_197 ),
	.I1(\top/processor/sha_core/n342_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n342_213 )
);
MUX2_LUT7 \top/processor/sha_core/n342_s191  (
	.I0(\top/processor/sha_core/n342_201 ),
	.I1(\top/processor/sha_core/n342_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n342_215 )
);
MUX2_LUT7 \top/processor/sha_core/n342_s192  (
	.I0(\top/processor/sha_core/n342_205 ),
	.I1(\top/processor/sha_core/n342_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n342_217 )
);
MUX2_LUT7 \top/processor/sha_core/n342_s193  (
	.I0(\top/processor/sha_core/n342_209 ),
	.I1(\top/processor/sha_core/n342_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n342_219 )
);
MUX2_LUT7 \top/processor/sha_core/n343_s190  (
	.I0(\top/processor/sha_core/n343_197 ),
	.I1(\top/processor/sha_core/n343_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n343_213 )
);
MUX2_LUT7 \top/processor/sha_core/n343_s191  (
	.I0(\top/processor/sha_core/n343_201 ),
	.I1(\top/processor/sha_core/n343_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n343_215 )
);
MUX2_LUT7 \top/processor/sha_core/n343_s192  (
	.I0(\top/processor/sha_core/n343_205 ),
	.I1(\top/processor/sha_core/n343_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n343_217 )
);
MUX2_LUT7 \top/processor/sha_core/n343_s193  (
	.I0(\top/processor/sha_core/n343_209 ),
	.I1(\top/processor/sha_core/n343_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n343_219 )
);
MUX2_LUT7 \top/processor/sha_core/n344_s190  (
	.I0(\top/processor/sha_core/n344_197 ),
	.I1(\top/processor/sha_core/n344_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n344_213 )
);
MUX2_LUT7 \top/processor/sha_core/n344_s191  (
	.I0(\top/processor/sha_core/n344_201 ),
	.I1(\top/processor/sha_core/n344_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n344_215 )
);
MUX2_LUT7 \top/processor/sha_core/n344_s192  (
	.I0(\top/processor/sha_core/n344_205 ),
	.I1(\top/processor/sha_core/n344_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n344_217 )
);
MUX2_LUT7 \top/processor/sha_core/n344_s193  (
	.I0(\top/processor/sha_core/n344_209 ),
	.I1(\top/processor/sha_core/n344_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n344_219 )
);
MUX2_LUT7 \top/processor/sha_core/n345_s190  (
	.I0(\top/processor/sha_core/n345_197 ),
	.I1(\top/processor/sha_core/n345_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n345_213 )
);
MUX2_LUT7 \top/processor/sha_core/n345_s191  (
	.I0(\top/processor/sha_core/n345_201 ),
	.I1(\top/processor/sha_core/n345_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n345_215 )
);
MUX2_LUT7 \top/processor/sha_core/n345_s192  (
	.I0(\top/processor/sha_core/n345_205 ),
	.I1(\top/processor/sha_core/n345_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n345_217 )
);
MUX2_LUT7 \top/processor/sha_core/n345_s193  (
	.I0(\top/processor/sha_core/n345_209 ),
	.I1(\top/processor/sha_core/n345_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n345_219 )
);
MUX2_LUT7 \top/processor/sha_core/n346_s190  (
	.I0(\top/processor/sha_core/n346_197 ),
	.I1(\top/processor/sha_core/n346_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n346_213 )
);
MUX2_LUT7 \top/processor/sha_core/n346_s191  (
	.I0(\top/processor/sha_core/n346_201 ),
	.I1(\top/processor/sha_core/n346_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n346_215 )
);
MUX2_LUT7 \top/processor/sha_core/n346_s192  (
	.I0(\top/processor/sha_core/n346_205 ),
	.I1(\top/processor/sha_core/n346_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n346_217 )
);
MUX2_LUT7 \top/processor/sha_core/n346_s193  (
	.I0(\top/processor/sha_core/n346_209 ),
	.I1(\top/processor/sha_core/n346_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n346_219 )
);
MUX2_LUT7 \top/processor/sha_core/n347_s190  (
	.I0(\top/processor/sha_core/n347_197 ),
	.I1(\top/processor/sha_core/n347_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n347_213 )
);
MUX2_LUT7 \top/processor/sha_core/n347_s191  (
	.I0(\top/processor/sha_core/n347_201 ),
	.I1(\top/processor/sha_core/n347_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n347_215 )
);
MUX2_LUT7 \top/processor/sha_core/n347_s192  (
	.I0(\top/processor/sha_core/n347_205 ),
	.I1(\top/processor/sha_core/n347_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n347_217 )
);
MUX2_LUT7 \top/processor/sha_core/n347_s193  (
	.I0(\top/processor/sha_core/n347_209 ),
	.I1(\top/processor/sha_core/n347_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n347_219 )
);
MUX2_LUT7 \top/processor/sha_core/n348_s190  (
	.I0(\top/processor/sha_core/n348_197 ),
	.I1(\top/processor/sha_core/n348_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n348_213 )
);
MUX2_LUT7 \top/processor/sha_core/n348_s191  (
	.I0(\top/processor/sha_core/n348_201 ),
	.I1(\top/processor/sha_core/n348_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n348_215 )
);
MUX2_LUT7 \top/processor/sha_core/n348_s192  (
	.I0(\top/processor/sha_core/n348_205 ),
	.I1(\top/processor/sha_core/n348_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n348_217 )
);
MUX2_LUT7 \top/processor/sha_core/n348_s193  (
	.I0(\top/processor/sha_core/n348_209 ),
	.I1(\top/processor/sha_core/n348_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n348_219 )
);
MUX2_LUT7 \top/processor/sha_core/n349_s190  (
	.I0(\top/processor/sha_core/n349_197 ),
	.I1(\top/processor/sha_core/n349_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n349_213 )
);
MUX2_LUT7 \top/processor/sha_core/n349_s191  (
	.I0(\top/processor/sha_core/n349_201 ),
	.I1(\top/processor/sha_core/n349_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n349_215 )
);
MUX2_LUT7 \top/processor/sha_core/n349_s192  (
	.I0(\top/processor/sha_core/n349_205 ),
	.I1(\top/processor/sha_core/n349_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n349_217 )
);
MUX2_LUT7 \top/processor/sha_core/n349_s193  (
	.I0(\top/processor/sha_core/n349_209 ),
	.I1(\top/processor/sha_core/n349_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n349_219 )
);
MUX2_LUT7 \top/processor/sha_core/n350_s190  (
	.I0(\top/processor/sha_core/n350_197 ),
	.I1(\top/processor/sha_core/n350_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n350_213 )
);
MUX2_LUT7 \top/processor/sha_core/n350_s191  (
	.I0(\top/processor/sha_core/n350_201 ),
	.I1(\top/processor/sha_core/n350_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n350_215 )
);
MUX2_LUT7 \top/processor/sha_core/n350_s192  (
	.I0(\top/processor/sha_core/n350_205 ),
	.I1(\top/processor/sha_core/n350_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n350_217 )
);
MUX2_LUT7 \top/processor/sha_core/n350_s193  (
	.I0(\top/processor/sha_core/n350_209 ),
	.I1(\top/processor/sha_core/n350_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n350_219 )
);
MUX2_LUT7 \top/processor/sha_core/n351_s190  (
	.I0(\top/processor/sha_core/n351_197 ),
	.I1(\top/processor/sha_core/n351_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n351_213 )
);
MUX2_LUT7 \top/processor/sha_core/n351_s191  (
	.I0(\top/processor/sha_core/n351_201 ),
	.I1(\top/processor/sha_core/n351_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n351_215 )
);
MUX2_LUT7 \top/processor/sha_core/n351_s192  (
	.I0(\top/processor/sha_core/n351_205 ),
	.I1(\top/processor/sha_core/n351_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n351_217 )
);
MUX2_LUT7 \top/processor/sha_core/n351_s193  (
	.I0(\top/processor/sha_core/n351_209 ),
	.I1(\top/processor/sha_core/n351_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n351_219 )
);
MUX2_LUT7 \top/processor/sha_core/n352_s190  (
	.I0(\top/processor/sha_core/n352_197 ),
	.I1(\top/processor/sha_core/n352_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n352_213 )
);
MUX2_LUT7 \top/processor/sha_core/n352_s191  (
	.I0(\top/processor/sha_core/n352_201 ),
	.I1(\top/processor/sha_core/n352_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n352_215 )
);
MUX2_LUT7 \top/processor/sha_core/n352_s192  (
	.I0(\top/processor/sha_core/n352_205 ),
	.I1(\top/processor/sha_core/n352_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n352_217 )
);
MUX2_LUT7 \top/processor/sha_core/n352_s193  (
	.I0(\top/processor/sha_core/n352_209 ),
	.I1(\top/processor/sha_core/n352_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n352_219 )
);
MUX2_LUT7 \top/processor/sha_core/n353_s190  (
	.I0(\top/processor/sha_core/n353_197 ),
	.I1(\top/processor/sha_core/n353_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n353_213 )
);
MUX2_LUT7 \top/processor/sha_core/n353_s191  (
	.I0(\top/processor/sha_core/n353_201 ),
	.I1(\top/processor/sha_core/n353_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n353_215 )
);
MUX2_LUT7 \top/processor/sha_core/n353_s192  (
	.I0(\top/processor/sha_core/n353_205 ),
	.I1(\top/processor/sha_core/n353_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n353_217 )
);
MUX2_LUT7 \top/processor/sha_core/n353_s193  (
	.I0(\top/processor/sha_core/n353_209 ),
	.I1(\top/processor/sha_core/n353_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n353_219 )
);
MUX2_LUT7 \top/processor/sha_core/n354_s190  (
	.I0(\top/processor/sha_core/n354_197 ),
	.I1(\top/processor/sha_core/n354_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n354_213 )
);
MUX2_LUT7 \top/processor/sha_core/n354_s191  (
	.I0(\top/processor/sha_core/n354_201 ),
	.I1(\top/processor/sha_core/n354_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n354_215 )
);
MUX2_LUT7 \top/processor/sha_core/n354_s192  (
	.I0(\top/processor/sha_core/n354_205 ),
	.I1(\top/processor/sha_core/n354_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n354_217 )
);
MUX2_LUT7 \top/processor/sha_core/n354_s193  (
	.I0(\top/processor/sha_core/n354_209 ),
	.I1(\top/processor/sha_core/n354_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n354_219 )
);
MUX2_LUT7 \top/processor/sha_core/n355_s190  (
	.I0(\top/processor/sha_core/n355_197 ),
	.I1(\top/processor/sha_core/n355_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n355_213 )
);
MUX2_LUT7 \top/processor/sha_core/n355_s191  (
	.I0(\top/processor/sha_core/n355_201 ),
	.I1(\top/processor/sha_core/n355_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n355_215 )
);
MUX2_LUT7 \top/processor/sha_core/n355_s192  (
	.I0(\top/processor/sha_core/n355_205 ),
	.I1(\top/processor/sha_core/n355_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n355_217 )
);
MUX2_LUT7 \top/processor/sha_core/n355_s193  (
	.I0(\top/processor/sha_core/n355_209 ),
	.I1(\top/processor/sha_core/n355_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n355_219 )
);
MUX2_LUT7 \top/processor/sha_core/n356_s190  (
	.I0(\top/processor/sha_core/n356_197 ),
	.I1(\top/processor/sha_core/n356_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n356_213 )
);
MUX2_LUT7 \top/processor/sha_core/n356_s191  (
	.I0(\top/processor/sha_core/n356_201 ),
	.I1(\top/processor/sha_core/n356_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n356_215 )
);
MUX2_LUT7 \top/processor/sha_core/n356_s192  (
	.I0(\top/processor/sha_core/n356_205 ),
	.I1(\top/processor/sha_core/n356_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n356_217 )
);
MUX2_LUT7 \top/processor/sha_core/n356_s193  (
	.I0(\top/processor/sha_core/n356_209 ),
	.I1(\top/processor/sha_core/n356_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n356_219 )
);
MUX2_LUT7 \top/processor/sha_core/n357_s190  (
	.I0(\top/processor/sha_core/n357_197 ),
	.I1(\top/processor/sha_core/n357_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n357_213 )
);
MUX2_LUT7 \top/processor/sha_core/n357_s191  (
	.I0(\top/processor/sha_core/n357_201 ),
	.I1(\top/processor/sha_core/n357_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n357_215 )
);
MUX2_LUT7 \top/processor/sha_core/n357_s192  (
	.I0(\top/processor/sha_core/n357_205 ),
	.I1(\top/processor/sha_core/n357_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n357_217 )
);
MUX2_LUT7 \top/processor/sha_core/n357_s193  (
	.I0(\top/processor/sha_core/n357_209 ),
	.I1(\top/processor/sha_core/n357_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n357_219 )
);
MUX2_LUT7 \top/processor/sha_core/n358_s190  (
	.I0(\top/processor/sha_core/n358_197 ),
	.I1(\top/processor/sha_core/n358_199 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n358_213 )
);
MUX2_LUT7 \top/processor/sha_core/n358_s191  (
	.I0(\top/processor/sha_core/n358_201 ),
	.I1(\top/processor/sha_core/n358_203 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n358_215 )
);
MUX2_LUT7 \top/processor/sha_core/n358_s192  (
	.I0(\top/processor/sha_core/n358_205 ),
	.I1(\top/processor/sha_core/n358_207 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n358_217 )
);
MUX2_LUT7 \top/processor/sha_core/n358_s193  (
	.I0(\top/processor/sha_core/n358_209 ),
	.I1(\top/processor/sha_core/n358_211 ),
	.S0(\top/processor/sha_core/t [3]),
	.O(\top/processor/sha_core/n358_219 )
);
MUX2_LUT7 \top/processor/sha_core/n3488_s173  (
	.I0(\top/processor/sha_core/n3488_189 ),
	.I1(\top/processor/sha_core/n3488_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3488_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3489_s173  (
	.I0(\top/processor/sha_core/n3489_189 ),
	.I1(\top/processor/sha_core/n3489_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3489_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3490_s173  (
	.I0(\top/processor/sha_core/n3490_189 ),
	.I1(\top/processor/sha_core/n3490_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3490_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3491_s173  (
	.I0(\top/processor/sha_core/n3491_189 ),
	.I1(\top/processor/sha_core/n3491_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3491_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3492_s173  (
	.I0(\top/processor/sha_core/n3492_189 ),
	.I1(\top/processor/sha_core/n3492_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3492_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3493_s173  (
	.I0(\top/processor/sha_core/n3493_189 ),
	.I1(\top/processor/sha_core/n3493_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3493_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3494_s173  (
	.I0(\top/processor/sha_core/n3494_190 ),
	.I1(\top/processor/sha_core/n3494_192 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3494_194 )
);
MUX2_LUT7 \top/processor/sha_core/n3495_s173  (
	.I0(\top/processor/sha_core/n3495_189 ),
	.I1(\top/processor/sha_core/n3495_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3495_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3496_s173  (
	.I0(\top/processor/sha_core/n3496_189 ),
	.I1(\top/processor/sha_core/n3496_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3496_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3497_s173  (
	.I0(\top/processor/sha_core/n3497_189 ),
	.I1(\top/processor/sha_core/n3497_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3497_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3498_s173  (
	.I0(\top/processor/sha_core/n3498_189 ),
	.I1(\top/processor/sha_core/n3498_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3498_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3499_s173  (
	.I0(\top/processor/sha_core/n3499_189 ),
	.I1(\top/processor/sha_core/n3499_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3499_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3500_s173  (
	.I0(\top/processor/sha_core/n3500_189 ),
	.I1(\top/processor/sha_core/n3500_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3500_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3501_s173  (
	.I0(\top/processor/sha_core/n3501_189 ),
	.I1(\top/processor/sha_core/n3501_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3501_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3502_s173  (
	.I0(\top/processor/sha_core/n3502_189 ),
	.I1(\top/processor/sha_core/n3502_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3502_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3503_s173  (
	.I0(\top/processor/sha_core/n3503_189 ),
	.I1(\top/processor/sha_core/n3503_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3503_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3504_s173  (
	.I0(\top/processor/sha_core/n3504_189 ),
	.I1(\top/processor/sha_core/n3504_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3504_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3505_s173  (
	.I0(\top/processor/sha_core/n3505_189 ),
	.I1(\top/processor/sha_core/n3505_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3505_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3506_s173  (
	.I0(\top/processor/sha_core/n3506_189 ),
	.I1(\top/processor/sha_core/n3506_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3506_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3507_s173  (
	.I0(\top/processor/sha_core/n3507_189 ),
	.I1(\top/processor/sha_core/n3507_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3507_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3508_s173  (
	.I0(\top/processor/sha_core/n3508_189 ),
	.I1(\top/processor/sha_core/n3508_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3508_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3509_s173  (
	.I0(\top/processor/sha_core/n3509_189 ),
	.I1(\top/processor/sha_core/n3509_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3509_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3511_s173  (
	.I0(\top/processor/sha_core/n3511_189 ),
	.I1(\top/processor/sha_core/n3511_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3511_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3512_s173  (
	.I0(\top/processor/sha_core/n3512_189 ),
	.I1(\top/processor/sha_core/n3512_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3512_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3513_s173  (
	.I0(\top/processor/sha_core/n3513_189 ),
	.I1(\top/processor/sha_core/n3513_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3513_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3514_s173  (
	.I0(\top/processor/sha_core/n3514_189 ),
	.I1(\top/processor/sha_core/n3514_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3514_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3515_s173  (
	.I0(\top/processor/sha_core/n3515_189 ),
	.I1(\top/processor/sha_core/n3515_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3515_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3516_s173  (
	.I0(\top/processor/sha_core/n3516_189 ),
	.I1(\top/processor/sha_core/n3516_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3516_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3517_s173  (
	.I0(\top/processor/sha_core/n3517_189 ),
	.I1(\top/processor/sha_core/n3517_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3517_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3518_s173  (
	.I0(\top/processor/sha_core/n3518_189 ),
	.I1(\top/processor/sha_core/n3518_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3518_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3519_s173  (
	.I0(\top/processor/sha_core/n3519_189 ),
	.I1(\top/processor/sha_core/n3519_191 ),
	.S0(\top/processor/sha_core/n3459_9 ),
	.O(\top/processor/sha_core/n3519_193 )
);
MUX2_LUT7 \top/processor/sha_core/n3860_s125  (
	.I0(\top/processor/sha_core/n3860_141 ),
	.I1(\top/processor/sha_core/n3860_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3860_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3861_s125  (
	.I0(\top/processor/sha_core/n3861_141 ),
	.I1(\top/processor/sha_core/n3861_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3861_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3862_s125  (
	.I0(\top/processor/sha_core/n3862_141 ),
	.I1(\top/processor/sha_core/n3862_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3862_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3863_s125  (
	.I0(\top/processor/sha_core/n3863_141 ),
	.I1(\top/processor/sha_core/n3863_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3863_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3864_s125  (
	.I0(\top/processor/sha_core/n3864_141 ),
	.I1(\top/processor/sha_core/n3864_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3864_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3865_s125  (
	.I0(\top/processor/sha_core/n3865_141 ),
	.I1(\top/processor/sha_core/n3865_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3865_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3866_s125  (
	.I0(\top/processor/sha_core/n3866_141 ),
	.I1(\top/processor/sha_core/n3866_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3866_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3867_s125  (
	.I0(\top/processor/sha_core/n3867_141 ),
	.I1(\top/processor/sha_core/n3867_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3867_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3868_s125  (
	.I0(\top/processor/sha_core/n3868_141 ),
	.I1(\top/processor/sha_core/n3868_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3868_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3869_s125  (
	.I0(\top/processor/sha_core/n3869_141 ),
	.I1(\top/processor/sha_core/n3869_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3869_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3870_s125  (
	.I0(\top/processor/sha_core/n3870_141 ),
	.I1(\top/processor/sha_core/n3870_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3870_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3871_s125  (
	.I0(\top/processor/sha_core/n3871_141 ),
	.I1(\top/processor/sha_core/n3871_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3871_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3872_s125  (
	.I0(\top/processor/sha_core/n3872_141 ),
	.I1(\top/processor/sha_core/n3872_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3872_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3873_s125  (
	.I0(\top/processor/sha_core/n3873_141 ),
	.I1(\top/processor/sha_core/n3873_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3873_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3874_s125  (
	.I0(\top/processor/sha_core/n3874_141 ),
	.I1(\top/processor/sha_core/n3874_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3874_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3875_s125  (
	.I0(\top/processor/sha_core/n3875_141 ),
	.I1(\top/processor/sha_core/n3875_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3875_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3876_s125  (
	.I0(\top/processor/sha_core/n3876_141 ),
	.I1(\top/processor/sha_core/n3876_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3876_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3877_s125  (
	.I0(\top/processor/sha_core/n3877_141 ),
	.I1(\top/processor/sha_core/n3877_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3877_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3878_s125  (
	.I0(\top/processor/sha_core/n3878_141 ),
	.I1(\top/processor/sha_core/n3878_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3878_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3879_s125  (
	.I0(\top/processor/sha_core/n3879_141 ),
	.I1(\top/processor/sha_core/n3879_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3879_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3880_s125  (
	.I0(\top/processor/sha_core/n3880_141 ),
	.I1(\top/processor/sha_core/n3880_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3880_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3881_s125  (
	.I0(\top/processor/sha_core/n3881_141 ),
	.I1(\top/processor/sha_core/n3881_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3881_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3882_s125  (
	.I0(\top/processor/sha_core/n3882_141 ),
	.I1(\top/processor/sha_core/n3882_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3882_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3883_s125  (
	.I0(\top/processor/sha_core/n3883_141 ),
	.I1(\top/processor/sha_core/n3883_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3883_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3884_s125  (
	.I0(\top/processor/sha_core/n3884_141 ),
	.I1(\top/processor/sha_core/n3884_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3884_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3885_s125  (
	.I0(\top/processor/sha_core/n3885_141 ),
	.I1(\top/processor/sha_core/n3885_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3885_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3886_s125  (
	.I0(\top/processor/sha_core/n3886_141 ),
	.I1(\top/processor/sha_core/n3886_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3886_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3887_s125  (
	.I0(\top/processor/sha_core/n3887_141 ),
	.I1(\top/processor/sha_core/n3887_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3887_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3888_s125  (
	.I0(\top/processor/sha_core/n3888_141 ),
	.I1(\top/processor/sha_core/n3888_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3888_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3889_s125  (
	.I0(\top/processor/sha_core/n3889_141 ),
	.I1(\top/processor/sha_core/n3889_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3889_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3890_s125  (
	.I0(\top/processor/sha_core/n3890_141 ),
	.I1(\top/processor/sha_core/n3890_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3890_145 )
);
MUX2_LUT7 \top/processor/sha_core/n3891_s125  (
	.I0(\top/processor/sha_core/n3891_141 ),
	.I1(\top/processor/sha_core/n3891_143 ),
	.S0(\top/processor/sha_core/n3834_9 ),
	.O(\top/processor/sha_core/n3891_145 )
);
MUX2_LUT8 \top/processor/sha_core/n327_s187  (
	.I0(\top/processor/sha_core/n327_213 ),
	.I1(\top/processor/sha_core/n327_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n327_221 )
);
MUX2_LUT8 \top/processor/sha_core/n327_s188  (
	.I0(\top/processor/sha_core/n327_217 ),
	.I1(\top/processor/sha_core/n327_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n327_223 )
);
MUX2_LUT8 \top/processor/sha_core/n328_s187  (
	.I0(\top/processor/sha_core/n328_213 ),
	.I1(\top/processor/sha_core/n328_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n328_221 )
);
MUX2_LUT8 \top/processor/sha_core/n328_s188  (
	.I0(\top/processor/sha_core/n328_217 ),
	.I1(\top/processor/sha_core/n328_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n328_223 )
);
MUX2_LUT8 \top/processor/sha_core/n329_s187  (
	.I0(\top/processor/sha_core/n329_213 ),
	.I1(\top/processor/sha_core/n329_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n329_221 )
);
MUX2_LUT8 \top/processor/sha_core/n329_s188  (
	.I0(\top/processor/sha_core/n329_217 ),
	.I1(\top/processor/sha_core/n329_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n329_223 )
);
MUX2_LUT8 \top/processor/sha_core/n330_s187  (
	.I0(\top/processor/sha_core/n330_213 ),
	.I1(\top/processor/sha_core/n330_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n330_221 )
);
MUX2_LUT8 \top/processor/sha_core/n330_s188  (
	.I0(\top/processor/sha_core/n330_217 ),
	.I1(\top/processor/sha_core/n330_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n330_223 )
);
MUX2_LUT8 \top/processor/sha_core/n331_s187  (
	.I0(\top/processor/sha_core/n331_213 ),
	.I1(\top/processor/sha_core/n331_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n331_221 )
);
MUX2_LUT8 \top/processor/sha_core/n331_s188  (
	.I0(\top/processor/sha_core/n331_217 ),
	.I1(\top/processor/sha_core/n331_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n331_223 )
);
MUX2_LUT8 \top/processor/sha_core/n332_s187  (
	.I0(\top/processor/sha_core/n332_213 ),
	.I1(\top/processor/sha_core/n332_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n332_221 )
);
MUX2_LUT8 \top/processor/sha_core/n332_s188  (
	.I0(\top/processor/sha_core/n332_217 ),
	.I1(\top/processor/sha_core/n332_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n332_223 )
);
MUX2_LUT8 \top/processor/sha_core/n333_s187  (
	.I0(\top/processor/sha_core/n333_213 ),
	.I1(\top/processor/sha_core/n333_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n333_221 )
);
MUX2_LUT8 \top/processor/sha_core/n333_s188  (
	.I0(\top/processor/sha_core/n333_217 ),
	.I1(\top/processor/sha_core/n333_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n333_223 )
);
MUX2_LUT8 \top/processor/sha_core/n334_s187  (
	.I0(\top/processor/sha_core/n334_213 ),
	.I1(\top/processor/sha_core/n334_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n334_221 )
);
MUX2_LUT8 \top/processor/sha_core/n334_s188  (
	.I0(\top/processor/sha_core/n334_217 ),
	.I1(\top/processor/sha_core/n334_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n334_223 )
);
MUX2_LUT8 \top/processor/sha_core/n335_s187  (
	.I0(\top/processor/sha_core/n335_213 ),
	.I1(\top/processor/sha_core/n335_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n335_221 )
);
MUX2_LUT8 \top/processor/sha_core/n335_s188  (
	.I0(\top/processor/sha_core/n335_217 ),
	.I1(\top/processor/sha_core/n335_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n335_223 )
);
MUX2_LUT8 \top/processor/sha_core/n336_s187  (
	.I0(\top/processor/sha_core/n336_213 ),
	.I1(\top/processor/sha_core/n336_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n336_221 )
);
MUX2_LUT8 \top/processor/sha_core/n336_s188  (
	.I0(\top/processor/sha_core/n336_217 ),
	.I1(\top/processor/sha_core/n336_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n336_223 )
);
MUX2_LUT8 \top/processor/sha_core/n337_s187  (
	.I0(\top/processor/sha_core/n337_213 ),
	.I1(\top/processor/sha_core/n337_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n337_221 )
);
MUX2_LUT8 \top/processor/sha_core/n337_s188  (
	.I0(\top/processor/sha_core/n337_217 ),
	.I1(\top/processor/sha_core/n337_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n337_223 )
);
MUX2_LUT8 \top/processor/sha_core/n338_s187  (
	.I0(\top/processor/sha_core/n338_213 ),
	.I1(\top/processor/sha_core/n338_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n338_221 )
);
MUX2_LUT8 \top/processor/sha_core/n338_s188  (
	.I0(\top/processor/sha_core/n338_217 ),
	.I1(\top/processor/sha_core/n338_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n338_223 )
);
MUX2_LUT8 \top/processor/sha_core/n339_s187  (
	.I0(\top/processor/sha_core/n339_213 ),
	.I1(\top/processor/sha_core/n339_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n339_221 )
);
MUX2_LUT8 \top/processor/sha_core/n339_s188  (
	.I0(\top/processor/sha_core/n339_217 ),
	.I1(\top/processor/sha_core/n339_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n339_223 )
);
MUX2_LUT8 \top/processor/sha_core/n340_s187  (
	.I0(\top/processor/sha_core/n340_213 ),
	.I1(\top/processor/sha_core/n340_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n340_221 )
);
MUX2_LUT8 \top/processor/sha_core/n340_s188  (
	.I0(\top/processor/sha_core/n340_217 ),
	.I1(\top/processor/sha_core/n340_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n340_223 )
);
MUX2_LUT8 \top/processor/sha_core/n341_s187  (
	.I0(\top/processor/sha_core/n341_213 ),
	.I1(\top/processor/sha_core/n341_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n341_221 )
);
MUX2_LUT8 \top/processor/sha_core/n341_s188  (
	.I0(\top/processor/sha_core/n341_217 ),
	.I1(\top/processor/sha_core/n341_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n341_223 )
);
MUX2_LUT8 \top/processor/sha_core/n342_s187  (
	.I0(\top/processor/sha_core/n342_213 ),
	.I1(\top/processor/sha_core/n342_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n342_221 )
);
MUX2_LUT8 \top/processor/sha_core/n342_s188  (
	.I0(\top/processor/sha_core/n342_217 ),
	.I1(\top/processor/sha_core/n342_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n342_223 )
);
MUX2_LUT8 \top/processor/sha_core/n343_s187  (
	.I0(\top/processor/sha_core/n343_213 ),
	.I1(\top/processor/sha_core/n343_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n343_221 )
);
MUX2_LUT8 \top/processor/sha_core/n343_s188  (
	.I0(\top/processor/sha_core/n343_217 ),
	.I1(\top/processor/sha_core/n343_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n343_223 )
);
MUX2_LUT8 \top/processor/sha_core/n344_s187  (
	.I0(\top/processor/sha_core/n344_213 ),
	.I1(\top/processor/sha_core/n344_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n344_221 )
);
MUX2_LUT8 \top/processor/sha_core/n344_s188  (
	.I0(\top/processor/sha_core/n344_217 ),
	.I1(\top/processor/sha_core/n344_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n344_223 )
);
MUX2_LUT8 \top/processor/sha_core/n345_s187  (
	.I0(\top/processor/sha_core/n345_213 ),
	.I1(\top/processor/sha_core/n345_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n345_221 )
);
MUX2_LUT8 \top/processor/sha_core/n345_s188  (
	.I0(\top/processor/sha_core/n345_217 ),
	.I1(\top/processor/sha_core/n345_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n345_223 )
);
MUX2_LUT8 \top/processor/sha_core/n346_s187  (
	.I0(\top/processor/sha_core/n346_213 ),
	.I1(\top/processor/sha_core/n346_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n346_221 )
);
MUX2_LUT8 \top/processor/sha_core/n346_s188  (
	.I0(\top/processor/sha_core/n346_217 ),
	.I1(\top/processor/sha_core/n346_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n346_223 )
);
MUX2_LUT8 \top/processor/sha_core/n347_s187  (
	.I0(\top/processor/sha_core/n347_213 ),
	.I1(\top/processor/sha_core/n347_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n347_221 )
);
MUX2_LUT8 \top/processor/sha_core/n347_s188  (
	.I0(\top/processor/sha_core/n347_217 ),
	.I1(\top/processor/sha_core/n347_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n347_223 )
);
MUX2_LUT8 \top/processor/sha_core/n348_s187  (
	.I0(\top/processor/sha_core/n348_213 ),
	.I1(\top/processor/sha_core/n348_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n348_221 )
);
MUX2_LUT8 \top/processor/sha_core/n348_s188  (
	.I0(\top/processor/sha_core/n348_217 ),
	.I1(\top/processor/sha_core/n348_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n348_223 )
);
MUX2_LUT8 \top/processor/sha_core/n349_s187  (
	.I0(\top/processor/sha_core/n349_213 ),
	.I1(\top/processor/sha_core/n349_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n349_221 )
);
MUX2_LUT8 \top/processor/sha_core/n349_s188  (
	.I0(\top/processor/sha_core/n349_217 ),
	.I1(\top/processor/sha_core/n349_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n349_223 )
);
MUX2_LUT8 \top/processor/sha_core/n350_s187  (
	.I0(\top/processor/sha_core/n350_213 ),
	.I1(\top/processor/sha_core/n350_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n350_221 )
);
MUX2_LUT8 \top/processor/sha_core/n350_s188  (
	.I0(\top/processor/sha_core/n350_217 ),
	.I1(\top/processor/sha_core/n350_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n350_223 )
);
MUX2_LUT8 \top/processor/sha_core/n351_s187  (
	.I0(\top/processor/sha_core/n351_213 ),
	.I1(\top/processor/sha_core/n351_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n351_221 )
);
MUX2_LUT8 \top/processor/sha_core/n351_s188  (
	.I0(\top/processor/sha_core/n351_217 ),
	.I1(\top/processor/sha_core/n351_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n351_223 )
);
MUX2_LUT8 \top/processor/sha_core/n352_s187  (
	.I0(\top/processor/sha_core/n352_213 ),
	.I1(\top/processor/sha_core/n352_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n352_221 )
);
MUX2_LUT8 \top/processor/sha_core/n352_s188  (
	.I0(\top/processor/sha_core/n352_217 ),
	.I1(\top/processor/sha_core/n352_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n352_223 )
);
MUX2_LUT8 \top/processor/sha_core/n353_s187  (
	.I0(\top/processor/sha_core/n353_213 ),
	.I1(\top/processor/sha_core/n353_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n353_221 )
);
MUX2_LUT8 \top/processor/sha_core/n353_s188  (
	.I0(\top/processor/sha_core/n353_217 ),
	.I1(\top/processor/sha_core/n353_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n353_223 )
);
MUX2_LUT8 \top/processor/sha_core/n354_s187  (
	.I0(\top/processor/sha_core/n354_213 ),
	.I1(\top/processor/sha_core/n354_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n354_221 )
);
MUX2_LUT8 \top/processor/sha_core/n354_s188  (
	.I0(\top/processor/sha_core/n354_217 ),
	.I1(\top/processor/sha_core/n354_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n354_223 )
);
MUX2_LUT8 \top/processor/sha_core/n355_s187  (
	.I0(\top/processor/sha_core/n355_213 ),
	.I1(\top/processor/sha_core/n355_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n355_221 )
);
MUX2_LUT8 \top/processor/sha_core/n355_s188  (
	.I0(\top/processor/sha_core/n355_217 ),
	.I1(\top/processor/sha_core/n355_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n355_223 )
);
MUX2_LUT8 \top/processor/sha_core/n356_s187  (
	.I0(\top/processor/sha_core/n356_213 ),
	.I1(\top/processor/sha_core/n356_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n356_221 )
);
MUX2_LUT8 \top/processor/sha_core/n356_s188  (
	.I0(\top/processor/sha_core/n356_217 ),
	.I1(\top/processor/sha_core/n356_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n356_223 )
);
MUX2_LUT8 \top/processor/sha_core/n357_s187  (
	.I0(\top/processor/sha_core/n357_213 ),
	.I1(\top/processor/sha_core/n357_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n357_221 )
);
MUX2_LUT8 \top/processor/sha_core/n357_s188  (
	.I0(\top/processor/sha_core/n357_217 ),
	.I1(\top/processor/sha_core/n357_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n357_223 )
);
MUX2_LUT8 \top/processor/sha_core/n358_s187  (
	.I0(\top/processor/sha_core/n358_213 ),
	.I1(\top/processor/sha_core/n358_215 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n358_221 )
);
MUX2_LUT8 \top/processor/sha_core/n358_s188  (
	.I0(\top/processor/sha_core/n358_217 ),
	.I1(\top/processor/sha_core/n358_219 ),
	.S0(\top/processor/sha_core/t [4]),
	.O(\top/processor/sha_core/n358_223 )
);
MUX2_LUT6 \top/processor/sha_core/n3607_s159  (
	.I0(\top/processor/sha_core/n3607_183 ),
	.I1(\top/processor/sha_core/n3607_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3607_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3607_s168  (
	.I0(\top/processor/sha_core/n3607_187 ),
	.I1(\top/processor/sha_core/n3607_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3607_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3607_s169  (
	.I0(\top/processor/sha_core/n3607_191 ),
	.I1(\top/processor/sha_core/n3607_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3607_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3608_s159  (
	.I0(\top/processor/sha_core/n3608_183 ),
	.I1(\top/processor/sha_core/n3608_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3608_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3608_s166  (
	.I0(\top/processor/sha_core/n3608_187 ),
	.I1(\top/processor/sha_core/n3608_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3608_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3608_s167  (
	.I0(\top/processor/sha_core/n3608_191 ),
	.I1(\top/processor/sha_core/n3608_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3608_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3609_s159  (
	.I0(\top/processor/sha_core/n3609_183 ),
	.I1(\top/processor/sha_core/n3609_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3609_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3609_s166  (
	.I0(\top/processor/sha_core/n3609_187 ),
	.I1(\top/processor/sha_core/n3609_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3609_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3609_s167  (
	.I0(\top/processor/sha_core/n3609_191 ),
	.I1(\top/processor/sha_core/n3609_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3609_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3610_s159  (
	.I0(\top/processor/sha_core/n3610_183 ),
	.I1(\top/processor/sha_core/n3610_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3610_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3610_s166  (
	.I0(\top/processor/sha_core/n3610_187 ),
	.I1(\top/processor/sha_core/n3610_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3610_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3610_s167  (
	.I0(\top/processor/sha_core/n3610_191 ),
	.I1(\top/processor/sha_core/n3610_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3610_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3611_s159  (
	.I0(\top/processor/sha_core/n3611_183 ),
	.I1(\top/processor/sha_core/n3611_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3611_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3611_s166  (
	.I0(\top/processor/sha_core/n3611_187 ),
	.I1(\top/processor/sha_core/n3611_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3611_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3611_s167  (
	.I0(\top/processor/sha_core/n3611_191 ),
	.I1(\top/processor/sha_core/n3611_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3611_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3612_s159  (
	.I0(\top/processor/sha_core/n3612_183 ),
	.I1(\top/processor/sha_core/n3612_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3612_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3612_s166  (
	.I0(\top/processor/sha_core/n3612_187 ),
	.I1(\top/processor/sha_core/n3612_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3612_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3612_s167  (
	.I0(\top/processor/sha_core/n3612_191 ),
	.I1(\top/processor/sha_core/n3612_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3612_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3613_s159  (
	.I0(\top/processor/sha_core/n3613_183 ),
	.I1(\top/processor/sha_core/n3613_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3613_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3613_s166  (
	.I0(\top/processor/sha_core/n3613_187 ),
	.I1(\top/processor/sha_core/n3613_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3613_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3613_s167  (
	.I0(\top/processor/sha_core/n3613_191 ),
	.I1(\top/processor/sha_core/n3613_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3613_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3614_s159  (
	.I0(\top/processor/sha_core/n3614_183 ),
	.I1(\top/processor/sha_core/n3614_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3614_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3614_s166  (
	.I0(\top/processor/sha_core/n3614_187 ),
	.I1(\top/processor/sha_core/n3614_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3614_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3614_s167  (
	.I0(\top/processor/sha_core/n3614_191 ),
	.I1(\top/processor/sha_core/n3614_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3614_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3615_s159  (
	.I0(\top/processor/sha_core/n3615_183 ),
	.I1(\top/processor/sha_core/n3615_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3615_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3615_s166  (
	.I0(\top/processor/sha_core/n3615_187 ),
	.I1(\top/processor/sha_core/n3615_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3615_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3615_s167  (
	.I0(\top/processor/sha_core/n3615_191 ),
	.I1(\top/processor/sha_core/n3615_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3615_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3616_s159  (
	.I0(\top/processor/sha_core/n3616_183 ),
	.I1(\top/processor/sha_core/n3616_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3616_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3616_s166  (
	.I0(\top/processor/sha_core/n3616_187 ),
	.I1(\top/processor/sha_core/n3616_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3616_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3616_s167  (
	.I0(\top/processor/sha_core/n3616_191 ),
	.I1(\top/processor/sha_core/n3616_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3616_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3617_s159  (
	.I0(\top/processor/sha_core/n3617_183 ),
	.I1(\top/processor/sha_core/n3617_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3617_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3617_s166  (
	.I0(\top/processor/sha_core/n3617_187 ),
	.I1(\top/processor/sha_core/n3617_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3617_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3617_s167  (
	.I0(\top/processor/sha_core/n3617_191 ),
	.I1(\top/processor/sha_core/n3617_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3617_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3618_s159  (
	.I0(\top/processor/sha_core/n3618_183 ),
	.I1(\top/processor/sha_core/n3618_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3618_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3618_s166  (
	.I0(\top/processor/sha_core/n3618_187 ),
	.I1(\top/processor/sha_core/n3618_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3618_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3618_s167  (
	.I0(\top/processor/sha_core/n3618_191 ),
	.I1(\top/processor/sha_core/n3618_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3618_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3619_s159  (
	.I0(\top/processor/sha_core/n3619_183 ),
	.I1(\top/processor/sha_core/n3619_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3619_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3619_s166  (
	.I0(\top/processor/sha_core/n3619_187 ),
	.I1(\top/processor/sha_core/n3619_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3619_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3619_s167  (
	.I0(\top/processor/sha_core/n3619_191 ),
	.I1(\top/processor/sha_core/n3619_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3619_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3620_s159  (
	.I0(\top/processor/sha_core/n3620_183 ),
	.I1(\top/processor/sha_core/n3620_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3620_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3620_s166  (
	.I0(\top/processor/sha_core/n3620_187 ),
	.I1(\top/processor/sha_core/n3620_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3620_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3620_s167  (
	.I0(\top/processor/sha_core/n3620_191 ),
	.I1(\top/processor/sha_core/n3620_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3620_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3621_s159  (
	.I0(\top/processor/sha_core/n3621_183 ),
	.I1(\top/processor/sha_core/n3621_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3621_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3621_s166  (
	.I0(\top/processor/sha_core/n3621_187 ),
	.I1(\top/processor/sha_core/n3621_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3621_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3621_s167  (
	.I0(\top/processor/sha_core/n3621_191 ),
	.I1(\top/processor/sha_core/n3621_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3621_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3622_s159  (
	.I0(\top/processor/sha_core/n3622_183 ),
	.I1(\top/processor/sha_core/n3622_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3622_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3622_s166  (
	.I0(\top/processor/sha_core/n3622_187 ),
	.I1(\top/processor/sha_core/n3622_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3622_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3622_s167  (
	.I0(\top/processor/sha_core/n3622_191 ),
	.I1(\top/processor/sha_core/n3622_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3622_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3623_s159  (
	.I0(\top/processor/sha_core/n3623_183 ),
	.I1(\top/processor/sha_core/n3623_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3623_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3623_s166  (
	.I0(\top/processor/sha_core/n3623_187 ),
	.I1(\top/processor/sha_core/n3623_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3623_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3623_s167  (
	.I0(\top/processor/sha_core/n3623_191 ),
	.I1(\top/processor/sha_core/n3623_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3623_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3624_s159  (
	.I0(\top/processor/sha_core/n3624_183 ),
	.I1(\top/processor/sha_core/n3624_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3624_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3624_s166  (
	.I0(\top/processor/sha_core/n3624_187 ),
	.I1(\top/processor/sha_core/n3624_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3624_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3624_s167  (
	.I0(\top/processor/sha_core/n3624_191 ),
	.I1(\top/processor/sha_core/n3624_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3624_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3625_s159  (
	.I0(\top/processor/sha_core/n3625_183 ),
	.I1(\top/processor/sha_core/n3625_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3625_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3625_s166  (
	.I0(\top/processor/sha_core/n3625_187 ),
	.I1(\top/processor/sha_core/n3625_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3625_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3625_s167  (
	.I0(\top/processor/sha_core/n3625_191 ),
	.I1(\top/processor/sha_core/n3625_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3625_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3626_s159  (
	.I0(\top/processor/sha_core/n3626_183 ),
	.I1(\top/processor/sha_core/n3626_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3626_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3626_s166  (
	.I0(\top/processor/sha_core/n3626_187 ),
	.I1(\top/processor/sha_core/n3626_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3626_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3626_s167  (
	.I0(\top/processor/sha_core/n3626_191 ),
	.I1(\top/processor/sha_core/n3626_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3626_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3627_s159  (
	.I0(\top/processor/sha_core/n3627_183 ),
	.I1(\top/processor/sha_core/n3627_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3627_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3627_s166  (
	.I0(\top/processor/sha_core/n3627_187 ),
	.I1(\top/processor/sha_core/n3627_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3627_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3627_s167  (
	.I0(\top/processor/sha_core/n3627_191 ),
	.I1(\top/processor/sha_core/n3627_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3627_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3628_s159  (
	.I0(\top/processor/sha_core/n3628_183 ),
	.I1(\top/processor/sha_core/n3628_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3628_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3628_s166  (
	.I0(\top/processor/sha_core/n3628_187 ),
	.I1(\top/processor/sha_core/n3628_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3628_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3628_s167  (
	.I0(\top/processor/sha_core/n3628_191 ),
	.I1(\top/processor/sha_core/n3628_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3628_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3629_s159  (
	.I0(\top/processor/sha_core/n3629_183 ),
	.I1(\top/processor/sha_core/n3629_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3629_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3629_s166  (
	.I0(\top/processor/sha_core/n3629_187 ),
	.I1(\top/processor/sha_core/n3629_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3629_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3629_s167  (
	.I0(\top/processor/sha_core/n3629_191 ),
	.I1(\top/processor/sha_core/n3629_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3629_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3630_s159  (
	.I0(\top/processor/sha_core/n3630_183 ),
	.I1(\top/processor/sha_core/n3630_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3630_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3630_s166  (
	.I0(\top/processor/sha_core/n3630_187 ),
	.I1(\top/processor/sha_core/n3630_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3630_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3630_s167  (
	.I0(\top/processor/sha_core/n3630_191 ),
	.I1(\top/processor/sha_core/n3630_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3630_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3631_s159  (
	.I0(\top/processor/sha_core/n3631_183 ),
	.I1(\top/processor/sha_core/n3631_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3631_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3631_s166  (
	.I0(\top/processor/sha_core/n3631_187 ),
	.I1(\top/processor/sha_core/n3631_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3631_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3631_s167  (
	.I0(\top/processor/sha_core/n3631_191 ),
	.I1(\top/processor/sha_core/n3631_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3631_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3632_s159  (
	.I0(\top/processor/sha_core/n3632_183 ),
	.I1(\top/processor/sha_core/n3632_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3632_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3632_s166  (
	.I0(\top/processor/sha_core/n3632_187 ),
	.I1(\top/processor/sha_core/n3632_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3632_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3632_s167  (
	.I0(\top/processor/sha_core/n3632_191 ),
	.I1(\top/processor/sha_core/n3632_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3632_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3633_s159  (
	.I0(\top/processor/sha_core/n3633_183 ),
	.I1(\top/processor/sha_core/n3633_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3633_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3633_s166  (
	.I0(\top/processor/sha_core/n3633_187 ),
	.I1(\top/processor/sha_core/n3633_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3633_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3633_s167  (
	.I0(\top/processor/sha_core/n3633_191 ),
	.I1(\top/processor/sha_core/n3633_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3633_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3634_s159  (
	.I0(\top/processor/sha_core/n3634_183 ),
	.I1(\top/processor/sha_core/n3634_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3634_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3634_s166  (
	.I0(\top/processor/sha_core/n3634_187 ),
	.I1(\top/processor/sha_core/n3634_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3634_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3634_s167  (
	.I0(\top/processor/sha_core/n3634_191 ),
	.I1(\top/processor/sha_core/n3634_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3634_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3635_s159  (
	.I0(\top/processor/sha_core/n3635_183 ),
	.I1(\top/processor/sha_core/n3635_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3635_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3635_s166  (
	.I0(\top/processor/sha_core/n3635_187 ),
	.I1(\top/processor/sha_core/n3635_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3635_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3635_s167  (
	.I0(\top/processor/sha_core/n3635_191 ),
	.I1(\top/processor/sha_core/n3635_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3635_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3636_s159  (
	.I0(\top/processor/sha_core/n3636_183 ),
	.I1(\top/processor/sha_core/n3636_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3636_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3636_s166  (
	.I0(\top/processor/sha_core/n3636_187 ),
	.I1(\top/processor/sha_core/n3636_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3636_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3636_s167  (
	.I0(\top/processor/sha_core/n3636_191 ),
	.I1(\top/processor/sha_core/n3636_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3636_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3637_s159  (
	.I0(\top/processor/sha_core/n3637_183 ),
	.I1(\top/processor/sha_core/n3637_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3637_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3637_s166  (
	.I0(\top/processor/sha_core/n3637_187 ),
	.I1(\top/processor/sha_core/n3637_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3637_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3637_s167  (
	.I0(\top/processor/sha_core/n3637_191 ),
	.I1(\top/processor/sha_core/n3637_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3637_185 )
);
MUX2_LUT6 \top/processor/sha_core/n3638_s159  (
	.I0(\top/processor/sha_core/n3638_183 ),
	.I1(\top/processor/sha_core/n3638_185 ),
	.S0(\top/processor/sha_core/n3577_11 ),
	.O(\top/processor/sha_core/n3638_181 )
);
MUX2_LUT5 \top/processor/sha_core/n3638_s166  (
	.I0(\top/processor/sha_core/n3638_187 ),
	.I1(\top/processor/sha_core/n3638_189 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3638_183 )
);
MUX2_LUT5 \top/processor/sha_core/n3638_s167  (
	.I0(\top/processor/sha_core/n3638_191 ),
	.I1(\top/processor/sha_core/n3638_193 ),
	.S0(\top/processor/sha_core/n3578_11 ),
	.O(\top/processor/sha_core/n3638_185 )
);
endmodule
